magic
tech sky130A
magscale 1 2
timestamp 1698659501
<< nwell >>
rect -3329 104 3425 142
rect -3425 -104 3425 104
rect -3425 -142 3329 -104
<< pmos >>
rect -3327 -42 -3297 42
rect -3231 -42 -3201 42
rect -3135 -42 -3105 42
rect -3039 -42 -3009 42
rect -2943 -42 -2913 42
rect -2847 -42 -2817 42
rect -2751 -42 -2721 42
rect -2655 -42 -2625 42
rect -2559 -42 -2529 42
rect -2463 -42 -2433 42
rect -2367 -42 -2337 42
rect -2271 -42 -2241 42
rect -2175 -42 -2145 42
rect -2079 -42 -2049 42
rect -1983 -42 -1953 42
rect -1887 -42 -1857 42
rect -1791 -42 -1761 42
rect -1695 -42 -1665 42
rect -1599 -42 -1569 42
rect -1503 -42 -1473 42
rect -1407 -42 -1377 42
rect -1311 -42 -1281 42
rect -1215 -42 -1185 42
rect -1119 -42 -1089 42
rect -1023 -42 -993 42
rect -927 -42 -897 42
rect -831 -42 -801 42
rect -735 -42 -705 42
rect -639 -42 -609 42
rect -543 -42 -513 42
rect -447 -42 -417 42
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
rect 417 -42 447 42
rect 513 -42 543 42
rect 609 -42 639 42
rect 705 -42 735 42
rect 801 -42 831 42
rect 897 -42 927 42
rect 993 -42 1023 42
rect 1089 -42 1119 42
rect 1185 -42 1215 42
rect 1281 -42 1311 42
rect 1377 -42 1407 42
rect 1473 -42 1503 42
rect 1569 -42 1599 42
rect 1665 -42 1695 42
rect 1761 -42 1791 42
rect 1857 -42 1887 42
rect 1953 -42 1983 42
rect 2049 -42 2079 42
rect 2145 -42 2175 42
rect 2241 -42 2271 42
rect 2337 -42 2367 42
rect 2433 -42 2463 42
rect 2529 -42 2559 42
rect 2625 -42 2655 42
rect 2721 -42 2751 42
rect 2817 -42 2847 42
rect 2913 -42 2943 42
rect 3009 -42 3039 42
rect 3105 -42 3135 42
rect 3201 -42 3231 42
rect 3297 -42 3327 42
<< pdiff >>
rect -3389 30 -3327 42
rect -3389 -30 -3377 30
rect -3343 -30 -3327 30
rect -3389 -42 -3327 -30
rect -3297 30 -3231 42
rect -3297 -30 -3281 30
rect -3247 -30 -3231 30
rect -3297 -42 -3231 -30
rect -3201 30 -3135 42
rect -3201 -30 -3185 30
rect -3151 -30 -3135 30
rect -3201 -42 -3135 -30
rect -3105 30 -3039 42
rect -3105 -30 -3089 30
rect -3055 -30 -3039 30
rect -3105 -42 -3039 -30
rect -3009 30 -2943 42
rect -3009 -30 -2993 30
rect -2959 -30 -2943 30
rect -3009 -42 -2943 -30
rect -2913 30 -2847 42
rect -2913 -30 -2897 30
rect -2863 -30 -2847 30
rect -2913 -42 -2847 -30
rect -2817 30 -2751 42
rect -2817 -30 -2801 30
rect -2767 -30 -2751 30
rect -2817 -42 -2751 -30
rect -2721 30 -2655 42
rect -2721 -30 -2705 30
rect -2671 -30 -2655 30
rect -2721 -42 -2655 -30
rect -2625 30 -2559 42
rect -2625 -30 -2609 30
rect -2575 -30 -2559 30
rect -2625 -42 -2559 -30
rect -2529 30 -2463 42
rect -2529 -30 -2513 30
rect -2479 -30 -2463 30
rect -2529 -42 -2463 -30
rect -2433 30 -2367 42
rect -2433 -30 -2417 30
rect -2383 -30 -2367 30
rect -2433 -42 -2367 -30
rect -2337 30 -2271 42
rect -2337 -30 -2321 30
rect -2287 -30 -2271 30
rect -2337 -42 -2271 -30
rect -2241 30 -2175 42
rect -2241 -30 -2225 30
rect -2191 -30 -2175 30
rect -2241 -42 -2175 -30
rect -2145 30 -2079 42
rect -2145 -30 -2129 30
rect -2095 -30 -2079 30
rect -2145 -42 -2079 -30
rect -2049 30 -1983 42
rect -2049 -30 -2033 30
rect -1999 -30 -1983 30
rect -2049 -42 -1983 -30
rect -1953 30 -1887 42
rect -1953 -30 -1937 30
rect -1903 -30 -1887 30
rect -1953 -42 -1887 -30
rect -1857 30 -1791 42
rect -1857 -30 -1841 30
rect -1807 -30 -1791 30
rect -1857 -42 -1791 -30
rect -1761 30 -1695 42
rect -1761 -30 -1745 30
rect -1711 -30 -1695 30
rect -1761 -42 -1695 -30
rect -1665 30 -1599 42
rect -1665 -30 -1649 30
rect -1615 -30 -1599 30
rect -1665 -42 -1599 -30
rect -1569 30 -1503 42
rect -1569 -30 -1553 30
rect -1519 -30 -1503 30
rect -1569 -42 -1503 -30
rect -1473 30 -1407 42
rect -1473 -30 -1457 30
rect -1423 -30 -1407 30
rect -1473 -42 -1407 -30
rect -1377 30 -1311 42
rect -1377 -30 -1361 30
rect -1327 -30 -1311 30
rect -1377 -42 -1311 -30
rect -1281 30 -1215 42
rect -1281 -30 -1265 30
rect -1231 -30 -1215 30
rect -1281 -42 -1215 -30
rect -1185 30 -1119 42
rect -1185 -30 -1169 30
rect -1135 -30 -1119 30
rect -1185 -42 -1119 -30
rect -1089 30 -1023 42
rect -1089 -30 -1073 30
rect -1039 -30 -1023 30
rect -1089 -42 -1023 -30
rect -993 30 -927 42
rect -993 -30 -977 30
rect -943 -30 -927 30
rect -993 -42 -927 -30
rect -897 30 -831 42
rect -897 -30 -881 30
rect -847 -30 -831 30
rect -897 -42 -831 -30
rect -801 30 -735 42
rect -801 -30 -785 30
rect -751 -30 -735 30
rect -801 -42 -735 -30
rect -705 30 -639 42
rect -705 -30 -689 30
rect -655 -30 -639 30
rect -705 -42 -639 -30
rect -609 30 -543 42
rect -609 -30 -593 30
rect -559 -30 -543 30
rect -609 -42 -543 -30
rect -513 30 -447 42
rect -513 -30 -497 30
rect -463 -30 -447 30
rect -513 -42 -447 -30
rect -417 30 -351 42
rect -417 -30 -401 30
rect -367 -30 -351 30
rect -417 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 417 42
rect 351 -30 367 30
rect 401 -30 417 30
rect 351 -42 417 -30
rect 447 30 513 42
rect 447 -30 463 30
rect 497 -30 513 30
rect 447 -42 513 -30
rect 543 30 609 42
rect 543 -30 559 30
rect 593 -30 609 30
rect 543 -42 609 -30
rect 639 30 705 42
rect 639 -30 655 30
rect 689 -30 705 30
rect 639 -42 705 -30
rect 735 30 801 42
rect 735 -30 751 30
rect 785 -30 801 30
rect 735 -42 801 -30
rect 831 30 897 42
rect 831 -30 847 30
rect 881 -30 897 30
rect 831 -42 897 -30
rect 927 30 993 42
rect 927 -30 943 30
rect 977 -30 993 30
rect 927 -42 993 -30
rect 1023 30 1089 42
rect 1023 -30 1039 30
rect 1073 -30 1089 30
rect 1023 -42 1089 -30
rect 1119 30 1185 42
rect 1119 -30 1135 30
rect 1169 -30 1185 30
rect 1119 -42 1185 -30
rect 1215 30 1281 42
rect 1215 -30 1231 30
rect 1265 -30 1281 30
rect 1215 -42 1281 -30
rect 1311 30 1377 42
rect 1311 -30 1327 30
rect 1361 -30 1377 30
rect 1311 -42 1377 -30
rect 1407 30 1473 42
rect 1407 -30 1423 30
rect 1457 -30 1473 30
rect 1407 -42 1473 -30
rect 1503 30 1569 42
rect 1503 -30 1519 30
rect 1553 -30 1569 30
rect 1503 -42 1569 -30
rect 1599 30 1665 42
rect 1599 -30 1615 30
rect 1649 -30 1665 30
rect 1599 -42 1665 -30
rect 1695 30 1761 42
rect 1695 -30 1711 30
rect 1745 -30 1761 30
rect 1695 -42 1761 -30
rect 1791 30 1857 42
rect 1791 -30 1807 30
rect 1841 -30 1857 30
rect 1791 -42 1857 -30
rect 1887 30 1953 42
rect 1887 -30 1903 30
rect 1937 -30 1953 30
rect 1887 -42 1953 -30
rect 1983 30 2049 42
rect 1983 -30 1999 30
rect 2033 -30 2049 30
rect 1983 -42 2049 -30
rect 2079 30 2145 42
rect 2079 -30 2095 30
rect 2129 -30 2145 30
rect 2079 -42 2145 -30
rect 2175 30 2241 42
rect 2175 -30 2191 30
rect 2225 -30 2241 30
rect 2175 -42 2241 -30
rect 2271 30 2337 42
rect 2271 -30 2287 30
rect 2321 -30 2337 30
rect 2271 -42 2337 -30
rect 2367 30 2433 42
rect 2367 -30 2383 30
rect 2417 -30 2433 30
rect 2367 -42 2433 -30
rect 2463 30 2529 42
rect 2463 -30 2479 30
rect 2513 -30 2529 30
rect 2463 -42 2529 -30
rect 2559 30 2625 42
rect 2559 -30 2575 30
rect 2609 -30 2625 30
rect 2559 -42 2625 -30
rect 2655 30 2721 42
rect 2655 -30 2671 30
rect 2705 -30 2721 30
rect 2655 -42 2721 -30
rect 2751 30 2817 42
rect 2751 -30 2767 30
rect 2801 -30 2817 30
rect 2751 -42 2817 -30
rect 2847 30 2913 42
rect 2847 -30 2863 30
rect 2897 -30 2913 30
rect 2847 -42 2913 -30
rect 2943 30 3009 42
rect 2943 -30 2959 30
rect 2993 -30 3009 30
rect 2943 -42 3009 -30
rect 3039 30 3105 42
rect 3039 -30 3055 30
rect 3089 -30 3105 30
rect 3039 -42 3105 -30
rect 3135 30 3201 42
rect 3135 -30 3151 30
rect 3185 -30 3201 30
rect 3135 -42 3201 -30
rect 3231 30 3297 42
rect 3231 -30 3247 30
rect 3281 -30 3297 30
rect 3231 -42 3297 -30
rect 3327 30 3389 42
rect 3327 -30 3343 30
rect 3377 -30 3389 30
rect 3327 -42 3389 -30
<< pdiffc >>
rect -3377 -30 -3343 30
rect -3281 -30 -3247 30
rect -3185 -30 -3151 30
rect -3089 -30 -3055 30
rect -2993 -30 -2959 30
rect -2897 -30 -2863 30
rect -2801 -30 -2767 30
rect -2705 -30 -2671 30
rect -2609 -30 -2575 30
rect -2513 -30 -2479 30
rect -2417 -30 -2383 30
rect -2321 -30 -2287 30
rect -2225 -30 -2191 30
rect -2129 -30 -2095 30
rect -2033 -30 -1999 30
rect -1937 -30 -1903 30
rect -1841 -30 -1807 30
rect -1745 -30 -1711 30
rect -1649 -30 -1615 30
rect -1553 -30 -1519 30
rect -1457 -30 -1423 30
rect -1361 -30 -1327 30
rect -1265 -30 -1231 30
rect -1169 -30 -1135 30
rect -1073 -30 -1039 30
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
rect 1039 -30 1073 30
rect 1135 -30 1169 30
rect 1231 -30 1265 30
rect 1327 -30 1361 30
rect 1423 -30 1457 30
rect 1519 -30 1553 30
rect 1615 -30 1649 30
rect 1711 -30 1745 30
rect 1807 -30 1841 30
rect 1903 -30 1937 30
rect 1999 -30 2033 30
rect 2095 -30 2129 30
rect 2191 -30 2225 30
rect 2287 -30 2321 30
rect 2383 -30 2417 30
rect 2479 -30 2513 30
rect 2575 -30 2609 30
rect 2671 -30 2705 30
rect 2767 -30 2801 30
rect 2863 -30 2897 30
rect 2959 -30 2993 30
rect 3055 -30 3089 30
rect 3151 -30 3185 30
rect 3247 -30 3281 30
rect 3343 -30 3377 30
<< poly >>
rect -3249 123 -3183 139
rect -3249 89 -3233 123
rect -3199 89 -3183 123
rect -3249 73 -3183 89
rect -3057 123 -2991 139
rect -3057 89 -3041 123
rect -3007 89 -2991 123
rect -3057 73 -2991 89
rect -2865 123 -2799 139
rect -2865 89 -2849 123
rect -2815 89 -2799 123
rect -2865 73 -2799 89
rect -2673 123 -2607 139
rect -2673 89 -2657 123
rect -2623 89 -2607 123
rect -2673 73 -2607 89
rect -2481 123 -2415 139
rect -2481 89 -2465 123
rect -2431 89 -2415 123
rect -2481 73 -2415 89
rect -2289 123 -2223 139
rect -2289 89 -2273 123
rect -2239 89 -2223 123
rect -2289 73 -2223 89
rect -2097 123 -2031 139
rect -2097 89 -2081 123
rect -2047 89 -2031 123
rect -2097 73 -2031 89
rect -1905 123 -1839 139
rect -1905 89 -1889 123
rect -1855 89 -1839 123
rect -1905 73 -1839 89
rect -1713 123 -1647 139
rect -1713 89 -1697 123
rect -1663 89 -1647 123
rect -1713 73 -1647 89
rect -1521 123 -1455 139
rect -1521 89 -1505 123
rect -1471 89 -1455 123
rect -1521 73 -1455 89
rect -1329 123 -1263 139
rect -1329 89 -1313 123
rect -1279 89 -1263 123
rect -1329 73 -1263 89
rect -1137 123 -1071 139
rect -1137 89 -1121 123
rect -1087 89 -1071 123
rect -1137 73 -1071 89
rect -945 123 -879 139
rect -945 89 -929 123
rect -895 89 -879 123
rect -945 73 -879 89
rect -753 123 -687 139
rect -753 89 -737 123
rect -703 89 -687 123
rect -753 73 -687 89
rect -561 123 -495 139
rect -561 89 -545 123
rect -511 89 -495 123
rect -561 73 -495 89
rect -369 123 -303 139
rect -369 89 -353 123
rect -319 89 -303 123
rect -369 73 -303 89
rect -177 123 -111 139
rect -177 89 -161 123
rect -127 89 -111 123
rect -177 73 -111 89
rect 15 123 81 139
rect 15 89 31 123
rect 65 89 81 123
rect 15 73 81 89
rect 207 123 273 139
rect 207 89 223 123
rect 257 89 273 123
rect 207 73 273 89
rect 399 123 465 139
rect 399 89 415 123
rect 449 89 465 123
rect 399 73 465 89
rect 591 123 657 139
rect 591 89 607 123
rect 641 89 657 123
rect 591 73 657 89
rect 783 123 849 139
rect 783 89 799 123
rect 833 89 849 123
rect 783 73 849 89
rect 975 123 1041 139
rect 975 89 991 123
rect 1025 89 1041 123
rect 975 73 1041 89
rect 1167 123 1233 139
rect 1167 89 1183 123
rect 1217 89 1233 123
rect 1167 73 1233 89
rect 1359 123 1425 139
rect 1359 89 1375 123
rect 1409 89 1425 123
rect 1359 73 1425 89
rect 1551 123 1617 139
rect 1551 89 1567 123
rect 1601 89 1617 123
rect 1551 73 1617 89
rect 1743 123 1809 139
rect 1743 89 1759 123
rect 1793 89 1809 123
rect 1743 73 1809 89
rect 1935 123 2001 139
rect 1935 89 1951 123
rect 1985 89 2001 123
rect 1935 73 2001 89
rect 2127 123 2193 139
rect 2127 89 2143 123
rect 2177 89 2193 123
rect 2127 73 2193 89
rect 2319 123 2385 139
rect 2319 89 2335 123
rect 2369 89 2385 123
rect 2319 73 2385 89
rect 2511 123 2577 139
rect 2511 89 2527 123
rect 2561 89 2577 123
rect 2511 73 2577 89
rect 2703 123 2769 139
rect 2703 89 2719 123
rect 2753 89 2769 123
rect 2703 73 2769 89
rect 2895 123 2961 139
rect 2895 89 2911 123
rect 2945 89 2961 123
rect 2895 73 2961 89
rect 3087 123 3153 139
rect 3087 89 3103 123
rect 3137 89 3153 123
rect 3087 73 3153 89
rect 3279 123 3345 139
rect 3279 89 3295 123
rect 3329 89 3345 123
rect 3279 73 3345 89
rect -3327 42 -3297 68
rect -3231 42 -3201 73
rect -3135 42 -3105 68
rect -3039 42 -3009 73
rect -2943 42 -2913 68
rect -2847 42 -2817 73
rect -2751 42 -2721 68
rect -2655 42 -2625 73
rect -2559 42 -2529 68
rect -2463 42 -2433 73
rect -2367 42 -2337 68
rect -2271 42 -2241 73
rect -2175 42 -2145 68
rect -2079 42 -2049 73
rect -1983 42 -1953 68
rect -1887 42 -1857 73
rect -1791 42 -1761 68
rect -1695 42 -1665 73
rect -1599 42 -1569 68
rect -1503 42 -1473 73
rect -1407 42 -1377 68
rect -1311 42 -1281 73
rect -1215 42 -1185 68
rect -1119 42 -1089 73
rect -1023 42 -993 68
rect -927 42 -897 73
rect -831 42 -801 68
rect -735 42 -705 73
rect -639 42 -609 68
rect -543 42 -513 73
rect -447 42 -417 68
rect -351 42 -321 73
rect -255 42 -225 68
rect -159 42 -129 73
rect -63 42 -33 68
rect 33 42 63 73
rect 129 42 159 68
rect 225 42 255 73
rect 321 42 351 68
rect 417 42 447 73
rect 513 42 543 68
rect 609 42 639 73
rect 705 42 735 68
rect 801 42 831 73
rect 897 42 927 68
rect 993 42 1023 73
rect 1089 42 1119 68
rect 1185 42 1215 73
rect 1281 42 1311 68
rect 1377 42 1407 73
rect 1473 42 1503 68
rect 1569 42 1599 73
rect 1665 42 1695 68
rect 1761 42 1791 73
rect 1857 42 1887 68
rect 1953 42 1983 73
rect 2049 42 2079 68
rect 2145 42 2175 73
rect 2241 42 2271 68
rect 2337 42 2367 73
rect 2433 42 2463 68
rect 2529 42 2559 73
rect 2625 42 2655 68
rect 2721 42 2751 73
rect 2817 42 2847 68
rect 2913 42 2943 73
rect 3009 42 3039 68
rect 3105 42 3135 73
rect 3201 42 3231 68
rect 3297 42 3327 73
rect -3327 -73 -3297 -42
rect -3231 -68 -3201 -42
rect -3135 -73 -3105 -42
rect -3039 -68 -3009 -42
rect -2943 -73 -2913 -42
rect -2847 -68 -2817 -42
rect -2751 -73 -2721 -42
rect -2655 -68 -2625 -42
rect -2559 -73 -2529 -42
rect -2463 -68 -2433 -42
rect -2367 -73 -2337 -42
rect -2271 -68 -2241 -42
rect -2175 -73 -2145 -42
rect -2079 -68 -2049 -42
rect -1983 -73 -1953 -42
rect -1887 -68 -1857 -42
rect -1791 -73 -1761 -42
rect -1695 -68 -1665 -42
rect -1599 -73 -1569 -42
rect -1503 -68 -1473 -42
rect -1407 -73 -1377 -42
rect -1311 -68 -1281 -42
rect -1215 -73 -1185 -42
rect -1119 -68 -1089 -42
rect -1023 -73 -993 -42
rect -927 -68 -897 -42
rect -831 -73 -801 -42
rect -735 -68 -705 -42
rect -639 -73 -609 -42
rect -543 -68 -513 -42
rect -447 -73 -417 -42
rect -351 -68 -321 -42
rect -255 -73 -225 -42
rect -159 -68 -129 -42
rect -63 -73 -33 -42
rect 33 -68 63 -42
rect 129 -73 159 -42
rect 225 -68 255 -42
rect 321 -73 351 -42
rect 417 -68 447 -42
rect 513 -73 543 -42
rect 609 -68 639 -42
rect 705 -73 735 -42
rect 801 -68 831 -42
rect 897 -73 927 -42
rect 993 -68 1023 -42
rect 1089 -73 1119 -42
rect 1185 -68 1215 -42
rect 1281 -73 1311 -42
rect 1377 -68 1407 -42
rect 1473 -73 1503 -42
rect 1569 -68 1599 -42
rect 1665 -73 1695 -42
rect 1761 -68 1791 -42
rect 1857 -73 1887 -42
rect 1953 -68 1983 -42
rect 2049 -73 2079 -42
rect 2145 -68 2175 -42
rect 2241 -73 2271 -42
rect 2337 -68 2367 -42
rect 2433 -73 2463 -42
rect 2529 -68 2559 -42
rect 2625 -73 2655 -42
rect 2721 -68 2751 -42
rect 2817 -73 2847 -42
rect 2913 -68 2943 -42
rect 3009 -73 3039 -42
rect 3105 -68 3135 -42
rect 3201 -73 3231 -42
rect 3297 -68 3327 -42
rect -3345 -89 -3279 -73
rect -3345 -123 -3329 -89
rect -3295 -123 -3279 -89
rect -3345 -139 -3279 -123
rect -3153 -89 -3087 -73
rect -3153 -123 -3137 -89
rect -3103 -123 -3087 -89
rect -3153 -139 -3087 -123
rect -2961 -89 -2895 -73
rect -2961 -123 -2945 -89
rect -2911 -123 -2895 -89
rect -2961 -139 -2895 -123
rect -2769 -89 -2703 -73
rect -2769 -123 -2753 -89
rect -2719 -123 -2703 -89
rect -2769 -139 -2703 -123
rect -2577 -89 -2511 -73
rect -2577 -123 -2561 -89
rect -2527 -123 -2511 -89
rect -2577 -139 -2511 -123
rect -2385 -89 -2319 -73
rect -2385 -123 -2369 -89
rect -2335 -123 -2319 -89
rect -2385 -139 -2319 -123
rect -2193 -89 -2127 -73
rect -2193 -123 -2177 -89
rect -2143 -123 -2127 -89
rect -2193 -139 -2127 -123
rect -2001 -89 -1935 -73
rect -2001 -123 -1985 -89
rect -1951 -123 -1935 -89
rect -2001 -139 -1935 -123
rect -1809 -89 -1743 -73
rect -1809 -123 -1793 -89
rect -1759 -123 -1743 -89
rect -1809 -139 -1743 -123
rect -1617 -89 -1551 -73
rect -1617 -123 -1601 -89
rect -1567 -123 -1551 -89
rect -1617 -139 -1551 -123
rect -1425 -89 -1359 -73
rect -1425 -123 -1409 -89
rect -1375 -123 -1359 -89
rect -1425 -139 -1359 -123
rect -1233 -89 -1167 -73
rect -1233 -123 -1217 -89
rect -1183 -123 -1167 -89
rect -1233 -139 -1167 -123
rect -1041 -89 -975 -73
rect -1041 -123 -1025 -89
rect -991 -123 -975 -89
rect -1041 -139 -975 -123
rect -849 -89 -783 -73
rect -849 -123 -833 -89
rect -799 -123 -783 -89
rect -849 -139 -783 -123
rect -657 -89 -591 -73
rect -657 -123 -641 -89
rect -607 -123 -591 -89
rect -657 -139 -591 -123
rect -465 -89 -399 -73
rect -465 -123 -449 -89
rect -415 -123 -399 -89
rect -465 -139 -399 -123
rect -273 -89 -207 -73
rect -273 -123 -257 -89
rect -223 -123 -207 -89
rect -273 -139 -207 -123
rect -81 -89 -15 -73
rect -81 -123 -65 -89
rect -31 -123 -15 -89
rect -81 -139 -15 -123
rect 111 -89 177 -73
rect 111 -123 127 -89
rect 161 -123 177 -89
rect 111 -139 177 -123
rect 303 -89 369 -73
rect 303 -123 319 -89
rect 353 -123 369 -89
rect 303 -139 369 -123
rect 495 -89 561 -73
rect 495 -123 511 -89
rect 545 -123 561 -89
rect 495 -139 561 -123
rect 687 -89 753 -73
rect 687 -123 703 -89
rect 737 -123 753 -89
rect 687 -139 753 -123
rect 879 -89 945 -73
rect 879 -123 895 -89
rect 929 -123 945 -89
rect 879 -139 945 -123
rect 1071 -89 1137 -73
rect 1071 -123 1087 -89
rect 1121 -123 1137 -89
rect 1071 -139 1137 -123
rect 1263 -89 1329 -73
rect 1263 -123 1279 -89
rect 1313 -123 1329 -89
rect 1263 -139 1329 -123
rect 1455 -89 1521 -73
rect 1455 -123 1471 -89
rect 1505 -123 1521 -89
rect 1455 -139 1521 -123
rect 1647 -89 1713 -73
rect 1647 -123 1663 -89
rect 1697 -123 1713 -89
rect 1647 -139 1713 -123
rect 1839 -89 1905 -73
rect 1839 -123 1855 -89
rect 1889 -123 1905 -89
rect 1839 -139 1905 -123
rect 2031 -89 2097 -73
rect 2031 -123 2047 -89
rect 2081 -123 2097 -89
rect 2031 -139 2097 -123
rect 2223 -89 2289 -73
rect 2223 -123 2239 -89
rect 2273 -123 2289 -89
rect 2223 -139 2289 -123
rect 2415 -89 2481 -73
rect 2415 -123 2431 -89
rect 2465 -123 2481 -89
rect 2415 -139 2481 -123
rect 2607 -89 2673 -73
rect 2607 -123 2623 -89
rect 2657 -123 2673 -89
rect 2607 -139 2673 -123
rect 2799 -89 2865 -73
rect 2799 -123 2815 -89
rect 2849 -123 2865 -89
rect 2799 -139 2865 -123
rect 2991 -89 3057 -73
rect 2991 -123 3007 -89
rect 3041 -123 3057 -89
rect 2991 -139 3057 -123
rect 3183 -89 3249 -73
rect 3183 -123 3199 -89
rect 3233 -123 3249 -89
rect 3183 -139 3249 -123
<< polycont >>
rect -3233 89 -3199 123
rect -3041 89 -3007 123
rect -2849 89 -2815 123
rect -2657 89 -2623 123
rect -2465 89 -2431 123
rect -2273 89 -2239 123
rect -2081 89 -2047 123
rect -1889 89 -1855 123
rect -1697 89 -1663 123
rect -1505 89 -1471 123
rect -1313 89 -1279 123
rect -1121 89 -1087 123
rect -929 89 -895 123
rect -737 89 -703 123
rect -545 89 -511 123
rect -353 89 -319 123
rect -161 89 -127 123
rect 31 89 65 123
rect 223 89 257 123
rect 415 89 449 123
rect 607 89 641 123
rect 799 89 833 123
rect 991 89 1025 123
rect 1183 89 1217 123
rect 1375 89 1409 123
rect 1567 89 1601 123
rect 1759 89 1793 123
rect 1951 89 1985 123
rect 2143 89 2177 123
rect 2335 89 2369 123
rect 2527 89 2561 123
rect 2719 89 2753 123
rect 2911 89 2945 123
rect 3103 89 3137 123
rect 3295 89 3329 123
rect -3329 -123 -3295 -89
rect -3137 -123 -3103 -89
rect -2945 -123 -2911 -89
rect -2753 -123 -2719 -89
rect -2561 -123 -2527 -89
rect -2369 -123 -2335 -89
rect -2177 -123 -2143 -89
rect -1985 -123 -1951 -89
rect -1793 -123 -1759 -89
rect -1601 -123 -1567 -89
rect -1409 -123 -1375 -89
rect -1217 -123 -1183 -89
rect -1025 -123 -991 -89
rect -833 -123 -799 -89
rect -641 -123 -607 -89
rect -449 -123 -415 -89
rect -257 -123 -223 -89
rect -65 -123 -31 -89
rect 127 -123 161 -89
rect 319 -123 353 -89
rect 511 -123 545 -89
rect 703 -123 737 -89
rect 895 -123 929 -89
rect 1087 -123 1121 -89
rect 1279 -123 1313 -89
rect 1471 -123 1505 -89
rect 1663 -123 1697 -89
rect 1855 -123 1889 -89
rect 2047 -123 2081 -89
rect 2239 -123 2273 -89
rect 2431 -123 2465 -89
rect 2623 -123 2657 -89
rect 2815 -123 2849 -89
rect 3007 -123 3041 -89
rect 3199 -123 3233 -89
<< locali >>
rect -3249 89 -3233 123
rect -3199 89 -3183 123
rect -3057 89 -3041 123
rect -3007 89 -2991 123
rect -2865 89 -2849 123
rect -2815 89 -2799 123
rect -2673 89 -2657 123
rect -2623 89 -2607 123
rect -2481 89 -2465 123
rect -2431 89 -2415 123
rect -2289 89 -2273 123
rect -2239 89 -2223 123
rect -2097 89 -2081 123
rect -2047 89 -2031 123
rect -1905 89 -1889 123
rect -1855 89 -1839 123
rect -1713 89 -1697 123
rect -1663 89 -1647 123
rect -1521 89 -1505 123
rect -1471 89 -1455 123
rect -1329 89 -1313 123
rect -1279 89 -1263 123
rect -1137 89 -1121 123
rect -1087 89 -1071 123
rect -945 89 -929 123
rect -895 89 -879 123
rect -753 89 -737 123
rect -703 89 -687 123
rect -561 89 -545 123
rect -511 89 -495 123
rect -369 89 -353 123
rect -319 89 -303 123
rect -177 89 -161 123
rect -127 89 -111 123
rect 15 89 31 123
rect 65 89 81 123
rect 207 89 223 123
rect 257 89 273 123
rect 399 89 415 123
rect 449 89 465 123
rect 591 89 607 123
rect 641 89 657 123
rect 783 89 799 123
rect 833 89 849 123
rect 975 89 991 123
rect 1025 89 1041 123
rect 1167 89 1183 123
rect 1217 89 1233 123
rect 1359 89 1375 123
rect 1409 89 1425 123
rect 1551 89 1567 123
rect 1601 89 1617 123
rect 1743 89 1759 123
rect 1793 89 1809 123
rect 1935 89 1951 123
rect 1985 89 2001 123
rect 2127 89 2143 123
rect 2177 89 2193 123
rect 2319 89 2335 123
rect 2369 89 2385 123
rect 2511 89 2527 123
rect 2561 89 2577 123
rect 2703 89 2719 123
rect 2753 89 2769 123
rect 2895 89 2911 123
rect 2945 89 2961 123
rect 3087 89 3103 123
rect 3137 89 3153 123
rect 3279 89 3295 123
rect 3329 89 3345 123
rect -3377 30 -3343 46
rect -3377 -46 -3343 -30
rect -3281 30 -3247 46
rect -3281 -46 -3247 -30
rect -3185 30 -3151 46
rect -3185 -46 -3151 -30
rect -3089 30 -3055 46
rect -3089 -46 -3055 -30
rect -2993 30 -2959 46
rect -2993 -46 -2959 -30
rect -2897 30 -2863 46
rect -2897 -46 -2863 -30
rect -2801 30 -2767 46
rect -2801 -46 -2767 -30
rect -2705 30 -2671 46
rect -2705 -46 -2671 -30
rect -2609 30 -2575 46
rect -2609 -46 -2575 -30
rect -2513 30 -2479 46
rect -2513 -46 -2479 -30
rect -2417 30 -2383 46
rect -2417 -46 -2383 -30
rect -2321 30 -2287 46
rect -2321 -46 -2287 -30
rect -2225 30 -2191 46
rect -2225 -46 -2191 -30
rect -2129 30 -2095 46
rect -2129 -46 -2095 -30
rect -2033 30 -1999 46
rect -2033 -46 -1999 -30
rect -1937 30 -1903 46
rect -1937 -46 -1903 -30
rect -1841 30 -1807 46
rect -1841 -46 -1807 -30
rect -1745 30 -1711 46
rect -1745 -46 -1711 -30
rect -1649 30 -1615 46
rect -1649 -46 -1615 -30
rect -1553 30 -1519 46
rect -1553 -46 -1519 -30
rect -1457 30 -1423 46
rect -1457 -46 -1423 -30
rect -1361 30 -1327 46
rect -1361 -46 -1327 -30
rect -1265 30 -1231 46
rect -1265 -46 -1231 -30
rect -1169 30 -1135 46
rect -1169 -46 -1135 -30
rect -1073 30 -1039 46
rect -1073 -46 -1039 -30
rect -977 30 -943 46
rect -977 -46 -943 -30
rect -881 30 -847 46
rect -881 -46 -847 -30
rect -785 30 -751 46
rect -785 -46 -751 -30
rect -689 30 -655 46
rect -689 -46 -655 -30
rect -593 30 -559 46
rect -593 -46 -559 -30
rect -497 30 -463 46
rect -497 -46 -463 -30
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect 463 30 497 46
rect 463 -46 497 -30
rect 559 30 593 46
rect 559 -46 593 -30
rect 655 30 689 46
rect 655 -46 689 -30
rect 751 30 785 46
rect 751 -46 785 -30
rect 847 30 881 46
rect 847 -46 881 -30
rect 943 30 977 46
rect 943 -46 977 -30
rect 1039 30 1073 46
rect 1039 -46 1073 -30
rect 1135 30 1169 46
rect 1135 -46 1169 -30
rect 1231 30 1265 46
rect 1231 -46 1265 -30
rect 1327 30 1361 46
rect 1327 -46 1361 -30
rect 1423 30 1457 46
rect 1423 -46 1457 -30
rect 1519 30 1553 46
rect 1519 -46 1553 -30
rect 1615 30 1649 46
rect 1615 -46 1649 -30
rect 1711 30 1745 46
rect 1711 -46 1745 -30
rect 1807 30 1841 46
rect 1807 -46 1841 -30
rect 1903 30 1937 46
rect 1903 -46 1937 -30
rect 1999 30 2033 46
rect 1999 -46 2033 -30
rect 2095 30 2129 46
rect 2095 -46 2129 -30
rect 2191 30 2225 46
rect 2191 -46 2225 -30
rect 2287 30 2321 46
rect 2287 -46 2321 -30
rect 2383 30 2417 46
rect 2383 -46 2417 -30
rect 2479 30 2513 46
rect 2479 -46 2513 -30
rect 2575 30 2609 46
rect 2575 -46 2609 -30
rect 2671 30 2705 46
rect 2671 -46 2705 -30
rect 2767 30 2801 46
rect 2767 -46 2801 -30
rect 2863 30 2897 46
rect 2863 -46 2897 -30
rect 2959 30 2993 46
rect 2959 -46 2993 -30
rect 3055 30 3089 46
rect 3055 -46 3089 -30
rect 3151 30 3185 46
rect 3151 -46 3185 -30
rect 3247 30 3281 46
rect 3247 -46 3281 -30
rect 3343 30 3377 46
rect 3343 -46 3377 -30
rect -3345 -123 -3329 -89
rect -3295 -123 -3279 -89
rect -3153 -123 -3137 -89
rect -3103 -123 -3087 -89
rect -2961 -123 -2945 -89
rect -2911 -123 -2895 -89
rect -2769 -123 -2753 -89
rect -2719 -123 -2703 -89
rect -2577 -123 -2561 -89
rect -2527 -123 -2511 -89
rect -2385 -123 -2369 -89
rect -2335 -123 -2319 -89
rect -2193 -123 -2177 -89
rect -2143 -123 -2127 -89
rect -2001 -123 -1985 -89
rect -1951 -123 -1935 -89
rect -1809 -123 -1793 -89
rect -1759 -123 -1743 -89
rect -1617 -123 -1601 -89
rect -1567 -123 -1551 -89
rect -1425 -123 -1409 -89
rect -1375 -123 -1359 -89
rect -1233 -123 -1217 -89
rect -1183 -123 -1167 -89
rect -1041 -123 -1025 -89
rect -991 -123 -975 -89
rect -849 -123 -833 -89
rect -799 -123 -783 -89
rect -657 -123 -641 -89
rect -607 -123 -591 -89
rect -465 -123 -449 -89
rect -415 -123 -399 -89
rect -273 -123 -257 -89
rect -223 -123 -207 -89
rect -81 -123 -65 -89
rect -31 -123 -15 -89
rect 111 -123 127 -89
rect 161 -123 177 -89
rect 303 -123 319 -89
rect 353 -123 369 -89
rect 495 -123 511 -89
rect 545 -123 561 -89
rect 687 -123 703 -89
rect 737 -123 753 -89
rect 879 -123 895 -89
rect 929 -123 945 -89
rect 1071 -123 1087 -89
rect 1121 -123 1137 -89
rect 1263 -123 1279 -89
rect 1313 -123 1329 -89
rect 1455 -123 1471 -89
rect 1505 -123 1521 -89
rect 1647 -123 1663 -89
rect 1697 -123 1713 -89
rect 1839 -123 1855 -89
rect 1889 -123 1905 -89
rect 2031 -123 2047 -89
rect 2081 -123 2097 -89
rect 2223 -123 2239 -89
rect 2273 -123 2289 -89
rect 2415 -123 2431 -89
rect 2465 -123 2481 -89
rect 2607 -123 2623 -89
rect 2657 -123 2673 -89
rect 2799 -123 2815 -89
rect 2849 -123 2865 -89
rect 2991 -123 3007 -89
rect 3041 -123 3057 -89
rect 3183 -123 3199 -89
rect 3233 -123 3249 -89
<< viali >>
rect -3377 -30 -3343 30
rect -3281 -30 -3247 30
rect -3185 -30 -3151 30
rect -3089 -30 -3055 30
rect -2993 -30 -2959 30
rect -2897 -30 -2863 30
rect -2801 -30 -2767 30
rect -2705 -30 -2671 30
rect -2609 -30 -2575 30
rect -2513 -30 -2479 30
rect -2417 -30 -2383 30
rect -2321 -30 -2287 30
rect -2225 -30 -2191 30
rect -2129 -30 -2095 30
rect -2033 -30 -1999 30
rect -1937 -30 -1903 30
rect -1841 -30 -1807 30
rect -1745 -30 -1711 30
rect -1649 -30 -1615 30
rect -1553 -30 -1519 30
rect -1457 -30 -1423 30
rect -1361 -30 -1327 30
rect -1265 -30 -1231 30
rect -1169 -30 -1135 30
rect -1073 -30 -1039 30
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
rect 1039 -30 1073 30
rect 1135 -30 1169 30
rect 1231 -30 1265 30
rect 1327 -30 1361 30
rect 1423 -30 1457 30
rect 1519 -30 1553 30
rect 1615 -30 1649 30
rect 1711 -30 1745 30
rect 1807 -30 1841 30
rect 1903 -30 1937 30
rect 1999 -30 2033 30
rect 2095 -30 2129 30
rect 2191 -30 2225 30
rect 2287 -30 2321 30
rect 2383 -30 2417 30
rect 2479 -30 2513 30
rect 2575 -30 2609 30
rect 2671 -30 2705 30
rect 2767 -30 2801 30
rect 2863 -30 2897 30
rect 2959 -30 2993 30
rect 3055 -30 3089 30
rect 3151 -30 3185 30
rect 3247 -30 3281 30
rect 3343 -30 3377 30
<< metal1 >>
rect -3383 30 -3337 42
rect -3383 -30 -3377 30
rect -3343 -30 -3337 30
rect -3383 -42 -3337 -30
rect -3287 30 -3241 42
rect -3287 -30 -3281 30
rect -3247 -30 -3241 30
rect -3287 -42 -3241 -30
rect -3191 30 -3145 42
rect -3191 -30 -3185 30
rect -3151 -30 -3145 30
rect -3191 -42 -3145 -30
rect -3095 30 -3049 42
rect -3095 -30 -3089 30
rect -3055 -30 -3049 30
rect -3095 -42 -3049 -30
rect -2999 30 -2953 42
rect -2999 -30 -2993 30
rect -2959 -30 -2953 30
rect -2999 -42 -2953 -30
rect -2903 30 -2857 42
rect -2903 -30 -2897 30
rect -2863 -30 -2857 30
rect -2903 -42 -2857 -30
rect -2807 30 -2761 42
rect -2807 -30 -2801 30
rect -2767 -30 -2761 30
rect -2807 -42 -2761 -30
rect -2711 30 -2665 42
rect -2711 -30 -2705 30
rect -2671 -30 -2665 30
rect -2711 -42 -2665 -30
rect -2615 30 -2569 42
rect -2615 -30 -2609 30
rect -2575 -30 -2569 30
rect -2615 -42 -2569 -30
rect -2519 30 -2473 42
rect -2519 -30 -2513 30
rect -2479 -30 -2473 30
rect -2519 -42 -2473 -30
rect -2423 30 -2377 42
rect -2423 -30 -2417 30
rect -2383 -30 -2377 30
rect -2423 -42 -2377 -30
rect -2327 30 -2281 42
rect -2327 -30 -2321 30
rect -2287 -30 -2281 30
rect -2327 -42 -2281 -30
rect -2231 30 -2185 42
rect -2231 -30 -2225 30
rect -2191 -30 -2185 30
rect -2231 -42 -2185 -30
rect -2135 30 -2089 42
rect -2135 -30 -2129 30
rect -2095 -30 -2089 30
rect -2135 -42 -2089 -30
rect -2039 30 -1993 42
rect -2039 -30 -2033 30
rect -1999 -30 -1993 30
rect -2039 -42 -1993 -30
rect -1943 30 -1897 42
rect -1943 -30 -1937 30
rect -1903 -30 -1897 30
rect -1943 -42 -1897 -30
rect -1847 30 -1801 42
rect -1847 -30 -1841 30
rect -1807 -30 -1801 30
rect -1847 -42 -1801 -30
rect -1751 30 -1705 42
rect -1751 -30 -1745 30
rect -1711 -30 -1705 30
rect -1751 -42 -1705 -30
rect -1655 30 -1609 42
rect -1655 -30 -1649 30
rect -1615 -30 -1609 30
rect -1655 -42 -1609 -30
rect -1559 30 -1513 42
rect -1559 -30 -1553 30
rect -1519 -30 -1513 30
rect -1559 -42 -1513 -30
rect -1463 30 -1417 42
rect -1463 -30 -1457 30
rect -1423 -30 -1417 30
rect -1463 -42 -1417 -30
rect -1367 30 -1321 42
rect -1367 -30 -1361 30
rect -1327 -30 -1321 30
rect -1367 -42 -1321 -30
rect -1271 30 -1225 42
rect -1271 -30 -1265 30
rect -1231 -30 -1225 30
rect -1271 -42 -1225 -30
rect -1175 30 -1129 42
rect -1175 -30 -1169 30
rect -1135 -30 -1129 30
rect -1175 -42 -1129 -30
rect -1079 30 -1033 42
rect -1079 -30 -1073 30
rect -1039 -30 -1033 30
rect -1079 -42 -1033 -30
rect -983 30 -937 42
rect -983 -30 -977 30
rect -943 -30 -937 30
rect -983 -42 -937 -30
rect -887 30 -841 42
rect -887 -30 -881 30
rect -847 -30 -841 30
rect -887 -42 -841 -30
rect -791 30 -745 42
rect -791 -30 -785 30
rect -751 -30 -745 30
rect -791 -42 -745 -30
rect -695 30 -649 42
rect -695 -30 -689 30
rect -655 -30 -649 30
rect -695 -42 -649 -30
rect -599 30 -553 42
rect -599 -30 -593 30
rect -559 -30 -553 30
rect -599 -42 -553 -30
rect -503 30 -457 42
rect -503 -30 -497 30
rect -463 -30 -457 30
rect -503 -42 -457 -30
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect 457 30 503 42
rect 457 -30 463 30
rect 497 -30 503 30
rect 457 -42 503 -30
rect 553 30 599 42
rect 553 -30 559 30
rect 593 -30 599 30
rect 553 -42 599 -30
rect 649 30 695 42
rect 649 -30 655 30
rect 689 -30 695 30
rect 649 -42 695 -30
rect 745 30 791 42
rect 745 -30 751 30
rect 785 -30 791 30
rect 745 -42 791 -30
rect 841 30 887 42
rect 841 -30 847 30
rect 881 -30 887 30
rect 841 -42 887 -30
rect 937 30 983 42
rect 937 -30 943 30
rect 977 -30 983 30
rect 937 -42 983 -30
rect 1033 30 1079 42
rect 1033 -30 1039 30
rect 1073 -30 1079 30
rect 1033 -42 1079 -30
rect 1129 30 1175 42
rect 1129 -30 1135 30
rect 1169 -30 1175 30
rect 1129 -42 1175 -30
rect 1225 30 1271 42
rect 1225 -30 1231 30
rect 1265 -30 1271 30
rect 1225 -42 1271 -30
rect 1321 30 1367 42
rect 1321 -30 1327 30
rect 1361 -30 1367 30
rect 1321 -42 1367 -30
rect 1417 30 1463 42
rect 1417 -30 1423 30
rect 1457 -30 1463 30
rect 1417 -42 1463 -30
rect 1513 30 1559 42
rect 1513 -30 1519 30
rect 1553 -30 1559 30
rect 1513 -42 1559 -30
rect 1609 30 1655 42
rect 1609 -30 1615 30
rect 1649 -30 1655 30
rect 1609 -42 1655 -30
rect 1705 30 1751 42
rect 1705 -30 1711 30
rect 1745 -30 1751 30
rect 1705 -42 1751 -30
rect 1801 30 1847 42
rect 1801 -30 1807 30
rect 1841 -30 1847 30
rect 1801 -42 1847 -30
rect 1897 30 1943 42
rect 1897 -30 1903 30
rect 1937 -30 1943 30
rect 1897 -42 1943 -30
rect 1993 30 2039 42
rect 1993 -30 1999 30
rect 2033 -30 2039 30
rect 1993 -42 2039 -30
rect 2089 30 2135 42
rect 2089 -30 2095 30
rect 2129 -30 2135 30
rect 2089 -42 2135 -30
rect 2185 30 2231 42
rect 2185 -30 2191 30
rect 2225 -30 2231 30
rect 2185 -42 2231 -30
rect 2281 30 2327 42
rect 2281 -30 2287 30
rect 2321 -30 2327 30
rect 2281 -42 2327 -30
rect 2377 30 2423 42
rect 2377 -30 2383 30
rect 2417 -30 2423 30
rect 2377 -42 2423 -30
rect 2473 30 2519 42
rect 2473 -30 2479 30
rect 2513 -30 2519 30
rect 2473 -42 2519 -30
rect 2569 30 2615 42
rect 2569 -30 2575 30
rect 2609 -30 2615 30
rect 2569 -42 2615 -30
rect 2665 30 2711 42
rect 2665 -30 2671 30
rect 2705 -30 2711 30
rect 2665 -42 2711 -30
rect 2761 30 2807 42
rect 2761 -30 2767 30
rect 2801 -30 2807 30
rect 2761 -42 2807 -30
rect 2857 30 2903 42
rect 2857 -30 2863 30
rect 2897 -30 2903 30
rect 2857 -42 2903 -30
rect 2953 30 2999 42
rect 2953 -30 2959 30
rect 2993 -30 2999 30
rect 2953 -42 2999 -30
rect 3049 30 3095 42
rect 3049 -30 3055 30
rect 3089 -30 3095 30
rect 3049 -42 3095 -30
rect 3145 30 3191 42
rect 3145 -30 3151 30
rect 3185 -30 3191 30
rect 3145 -42 3191 -30
rect 3241 30 3287 42
rect 3241 -30 3247 30
rect 3281 -30 3287 30
rect 3241 -42 3287 -30
rect 3337 30 3383 42
rect 3337 -30 3343 30
rect 3377 -30 3383 30
rect 3337 -42 3383 -30
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 70 diffcov 100 polycov 100 guard 0 glc 0 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
