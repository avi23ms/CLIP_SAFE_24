magic
tech sky130A
magscale 1 2
timestamp 1727642364
<< viali >>
rect 1944 306 1978 340
rect 114 216 148 250
rect 452 216 488 252
<< metal1 >>
rect 48 568 76 586
rect 1928 344 2004 350
rect 1928 340 2060 344
rect 1928 306 1944 340
rect 1978 306 2060 340
rect 1928 294 2060 306
rect 94 254 172 256
rect -147 250 172 254
rect -147 216 114 250
rect 148 216 172 250
rect 94 208 172 216
rect 438 252 504 262
rect 438 216 452 252
rect 488 216 504 252
rect 438 210 504 216
rect 452 170 488 210
rect -110 134 488 170
rect 28 -46 76 -16
use sky130_fd_sc_hd__xnor2_4  sky130_fd_sc_hd__xnor2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 0 0 1 0
box -38 -48 2062 592
<< labels >>
rlabel metal1 -116 236 -116 236 1 B
port 1 n
rlabel metal1 -104 158 -104 158 1 A
port 2 n
rlabel metal1 48 -32 48 -32 1 gnd
port 3 n
rlabel metal1 58 570 58 570 1 Vdd
port 4 n
<< end >>
