magic
tech sky130A
magscale 1 2
timestamp 1699103691
<< nwell >>
rect -1265 188 1265 226
rect -1361 -226 1361 188
<< pmos >>
rect -1263 -126 -1233 126
rect -1167 -126 -1137 126
rect -1071 -126 -1041 126
rect -975 -126 -945 126
rect -879 -126 -849 126
rect -783 -126 -753 126
rect -687 -126 -657 126
rect -591 -126 -561 126
rect -495 -126 -465 126
rect -399 -126 -369 126
rect -303 -126 -273 126
rect -207 -126 -177 126
rect -111 -126 -81 126
rect -15 -126 15 126
rect 81 -126 111 126
rect 177 -126 207 126
rect 273 -126 303 126
rect 369 -126 399 126
rect 465 -126 495 126
rect 561 -126 591 126
rect 657 -126 687 126
rect 753 -126 783 126
rect 849 -126 879 126
rect 945 -126 975 126
rect 1041 -126 1071 126
rect 1137 -126 1167 126
rect 1233 -126 1263 126
<< pdiff >>
rect -1325 114 -1263 126
rect -1325 -114 -1313 114
rect -1279 -114 -1263 114
rect -1325 -126 -1263 -114
rect -1233 114 -1167 126
rect -1233 -114 -1217 114
rect -1183 -114 -1167 114
rect -1233 -126 -1167 -114
rect -1137 114 -1071 126
rect -1137 -114 -1121 114
rect -1087 -114 -1071 114
rect -1137 -126 -1071 -114
rect -1041 114 -975 126
rect -1041 -114 -1025 114
rect -991 -114 -975 114
rect -1041 -126 -975 -114
rect -945 114 -879 126
rect -945 -114 -929 114
rect -895 -114 -879 114
rect -945 -126 -879 -114
rect -849 114 -783 126
rect -849 -114 -833 114
rect -799 -114 -783 114
rect -849 -126 -783 -114
rect -753 114 -687 126
rect -753 -114 -737 114
rect -703 -114 -687 114
rect -753 -126 -687 -114
rect -657 114 -591 126
rect -657 -114 -641 114
rect -607 -114 -591 114
rect -657 -126 -591 -114
rect -561 114 -495 126
rect -561 -114 -545 114
rect -511 -114 -495 114
rect -561 -126 -495 -114
rect -465 114 -399 126
rect -465 -114 -449 114
rect -415 -114 -399 114
rect -465 -126 -399 -114
rect -369 114 -303 126
rect -369 -114 -353 114
rect -319 -114 -303 114
rect -369 -126 -303 -114
rect -273 114 -207 126
rect -273 -114 -257 114
rect -223 -114 -207 114
rect -273 -126 -207 -114
rect -177 114 -111 126
rect -177 -114 -161 114
rect -127 -114 -111 114
rect -177 -126 -111 -114
rect -81 114 -15 126
rect -81 -114 -65 114
rect -31 -114 -15 114
rect -81 -126 -15 -114
rect 15 114 81 126
rect 15 -114 31 114
rect 65 -114 81 114
rect 15 -126 81 -114
rect 111 114 177 126
rect 111 -114 127 114
rect 161 -114 177 114
rect 111 -126 177 -114
rect 207 114 273 126
rect 207 -114 223 114
rect 257 -114 273 114
rect 207 -126 273 -114
rect 303 114 369 126
rect 303 -114 319 114
rect 353 -114 369 114
rect 303 -126 369 -114
rect 399 114 465 126
rect 399 -114 415 114
rect 449 -114 465 114
rect 399 -126 465 -114
rect 495 114 561 126
rect 495 -114 511 114
rect 545 -114 561 114
rect 495 -126 561 -114
rect 591 114 657 126
rect 591 -114 607 114
rect 641 -114 657 114
rect 591 -126 657 -114
rect 687 114 753 126
rect 687 -114 703 114
rect 737 -114 753 114
rect 687 -126 753 -114
rect 783 114 849 126
rect 783 -114 799 114
rect 833 -114 849 114
rect 783 -126 849 -114
rect 879 114 945 126
rect 879 -114 895 114
rect 929 -114 945 114
rect 879 -126 945 -114
rect 975 114 1041 126
rect 975 -114 991 114
rect 1025 -114 1041 114
rect 975 -126 1041 -114
rect 1071 114 1137 126
rect 1071 -114 1087 114
rect 1121 -114 1137 114
rect 1071 -126 1137 -114
rect 1167 114 1233 126
rect 1167 -114 1183 114
rect 1217 -114 1233 114
rect 1167 -126 1233 -114
rect 1263 114 1325 126
rect 1263 -114 1279 114
rect 1313 -114 1325 114
rect 1263 -126 1325 -114
<< pdiffc >>
rect -1313 -114 -1279 114
rect -1217 -114 -1183 114
rect -1121 -114 -1087 114
rect -1025 -114 -991 114
rect -929 -114 -895 114
rect -833 -114 -799 114
rect -737 -114 -703 114
rect -641 -114 -607 114
rect -545 -114 -511 114
rect -449 -114 -415 114
rect -353 -114 -319 114
rect -257 -114 -223 114
rect -161 -114 -127 114
rect -65 -114 -31 114
rect 31 -114 65 114
rect 127 -114 161 114
rect 223 -114 257 114
rect 319 -114 353 114
rect 415 -114 449 114
rect 511 -114 545 114
rect 607 -114 641 114
rect 703 -114 737 114
rect 799 -114 833 114
rect 895 -114 929 114
rect 991 -114 1025 114
rect 1087 -114 1121 114
rect 1183 -114 1217 114
rect 1279 -114 1313 114
<< poly >>
rect -1185 207 -1119 223
rect -1185 173 -1169 207
rect -1135 173 -1119 207
rect -1185 157 -1119 173
rect -993 207 -927 223
rect -993 173 -977 207
rect -943 173 -927 207
rect -993 157 -927 173
rect -801 207 -735 223
rect -801 173 -785 207
rect -751 173 -735 207
rect -801 157 -735 173
rect -609 207 -543 223
rect -609 173 -593 207
rect -559 173 -543 207
rect -609 157 -543 173
rect -417 207 -351 223
rect -417 173 -401 207
rect -367 173 -351 207
rect -417 157 -351 173
rect -225 207 -159 223
rect -225 173 -209 207
rect -175 173 -159 207
rect -225 157 -159 173
rect -33 207 33 223
rect -33 173 -17 207
rect 17 173 33 207
rect -33 157 33 173
rect 159 207 225 223
rect 159 173 175 207
rect 209 173 225 207
rect 159 157 225 173
rect 351 207 417 223
rect 351 173 367 207
rect 401 173 417 207
rect 351 157 417 173
rect 543 207 609 223
rect 543 173 559 207
rect 593 173 609 207
rect 543 157 609 173
rect 735 207 801 223
rect 735 173 751 207
rect 785 173 801 207
rect 735 157 801 173
rect 927 207 993 223
rect 927 173 943 207
rect 977 173 993 207
rect 927 157 993 173
rect 1119 207 1185 223
rect 1119 173 1135 207
rect 1169 173 1185 207
rect 1119 157 1185 173
rect -1263 126 -1233 152
rect -1167 126 -1137 157
rect -1071 126 -1041 152
rect -975 126 -945 157
rect -879 126 -849 152
rect -783 126 -753 157
rect -687 126 -657 152
rect -591 126 -561 157
rect -495 126 -465 152
rect -399 126 -369 157
rect -303 126 -273 152
rect -207 126 -177 157
rect -111 126 -81 152
rect -15 126 15 157
rect 81 126 111 152
rect 177 126 207 157
rect 273 126 303 152
rect 369 126 399 157
rect 465 126 495 152
rect 561 126 591 157
rect 657 126 687 152
rect 753 126 783 157
rect 849 126 879 152
rect 945 126 975 157
rect 1041 126 1071 152
rect 1137 126 1167 157
rect 1233 126 1263 152
rect -1263 -157 -1233 -126
rect -1167 -152 -1137 -126
rect -1071 -157 -1041 -126
rect -975 -152 -945 -126
rect -879 -157 -849 -126
rect -783 -152 -753 -126
rect -687 -157 -657 -126
rect -591 -152 -561 -126
rect -495 -157 -465 -126
rect -399 -152 -369 -126
rect -303 -157 -273 -126
rect -207 -152 -177 -126
rect -111 -157 -81 -126
rect -15 -152 15 -126
rect 81 -157 111 -126
rect 177 -152 207 -126
rect 273 -157 303 -126
rect 369 -152 399 -126
rect 465 -157 495 -126
rect 561 -152 591 -126
rect 657 -157 687 -126
rect 753 -152 783 -126
rect 849 -157 879 -126
rect 945 -152 975 -126
rect 1041 -157 1071 -126
rect 1137 -152 1167 -126
rect 1233 -157 1263 -126
rect -1281 -173 -1215 -157
rect -1281 -207 -1265 -173
rect -1231 -207 -1215 -173
rect -1281 -223 -1215 -207
rect -1089 -173 -1023 -157
rect -1089 -207 -1073 -173
rect -1039 -207 -1023 -173
rect -1089 -223 -1023 -207
rect -897 -173 -831 -157
rect -897 -207 -881 -173
rect -847 -207 -831 -173
rect -897 -223 -831 -207
rect -705 -173 -639 -157
rect -705 -207 -689 -173
rect -655 -207 -639 -173
rect -705 -223 -639 -207
rect -513 -173 -447 -157
rect -513 -207 -497 -173
rect -463 -207 -447 -173
rect -513 -223 -447 -207
rect -321 -173 -255 -157
rect -321 -207 -305 -173
rect -271 -207 -255 -173
rect -321 -223 -255 -207
rect -129 -173 -63 -157
rect -129 -207 -113 -173
rect -79 -207 -63 -173
rect -129 -223 -63 -207
rect 63 -173 129 -157
rect 63 -207 79 -173
rect 113 -207 129 -173
rect 63 -223 129 -207
rect 255 -173 321 -157
rect 255 -207 271 -173
rect 305 -207 321 -173
rect 255 -223 321 -207
rect 447 -173 513 -157
rect 447 -207 463 -173
rect 497 -207 513 -173
rect 447 -223 513 -207
rect 639 -173 705 -157
rect 639 -207 655 -173
rect 689 -207 705 -173
rect 639 -223 705 -207
rect 831 -173 897 -157
rect 831 -207 847 -173
rect 881 -207 897 -173
rect 831 -223 897 -207
rect 1023 -173 1089 -157
rect 1023 -207 1039 -173
rect 1073 -207 1089 -173
rect 1023 -223 1089 -207
rect 1215 -173 1281 -157
rect 1215 -207 1231 -173
rect 1265 -207 1281 -173
rect 1215 -223 1281 -207
<< polycont >>
rect -1169 173 -1135 207
rect -977 173 -943 207
rect -785 173 -751 207
rect -593 173 -559 207
rect -401 173 -367 207
rect -209 173 -175 207
rect -17 173 17 207
rect 175 173 209 207
rect 367 173 401 207
rect 559 173 593 207
rect 751 173 785 207
rect 943 173 977 207
rect 1135 173 1169 207
rect -1265 -207 -1231 -173
rect -1073 -207 -1039 -173
rect -881 -207 -847 -173
rect -689 -207 -655 -173
rect -497 -207 -463 -173
rect -305 -207 -271 -173
rect -113 -207 -79 -173
rect 79 -207 113 -173
rect 271 -207 305 -173
rect 463 -207 497 -173
rect 655 -207 689 -173
rect 847 -207 881 -173
rect 1039 -207 1073 -173
rect 1231 -207 1265 -173
<< locali >>
rect -1185 173 -1169 207
rect -1135 173 -1119 207
rect -993 173 -977 207
rect -943 173 -927 207
rect -801 173 -785 207
rect -751 173 -735 207
rect -609 173 -593 207
rect -559 173 -543 207
rect -417 173 -401 207
rect -367 173 -351 207
rect -225 173 -209 207
rect -175 173 -159 207
rect -33 173 -17 207
rect 17 173 33 207
rect 159 173 175 207
rect 209 173 225 207
rect 351 173 367 207
rect 401 173 417 207
rect 543 173 559 207
rect 593 173 609 207
rect 735 173 751 207
rect 785 173 801 207
rect 927 173 943 207
rect 977 173 993 207
rect 1119 173 1135 207
rect 1169 173 1185 207
rect -1313 114 -1279 130
rect -1313 -130 -1279 -114
rect -1217 114 -1183 130
rect -1217 -130 -1183 -114
rect -1121 114 -1087 130
rect -1121 -130 -1087 -114
rect -1025 114 -991 130
rect -1025 -130 -991 -114
rect -929 114 -895 130
rect -929 -130 -895 -114
rect -833 114 -799 130
rect -833 -130 -799 -114
rect -737 114 -703 130
rect -737 -130 -703 -114
rect -641 114 -607 130
rect -641 -130 -607 -114
rect -545 114 -511 130
rect -545 -130 -511 -114
rect -449 114 -415 130
rect -449 -130 -415 -114
rect -353 114 -319 130
rect -353 -130 -319 -114
rect -257 114 -223 130
rect -257 -130 -223 -114
rect -161 114 -127 130
rect -161 -130 -127 -114
rect -65 114 -31 130
rect -65 -130 -31 -114
rect 31 114 65 130
rect 31 -130 65 -114
rect 127 114 161 130
rect 127 -130 161 -114
rect 223 114 257 130
rect 223 -130 257 -114
rect 319 114 353 130
rect 319 -130 353 -114
rect 415 114 449 130
rect 415 -130 449 -114
rect 511 114 545 130
rect 511 -130 545 -114
rect 607 114 641 130
rect 607 -130 641 -114
rect 703 114 737 130
rect 703 -130 737 -114
rect 799 114 833 130
rect 799 -130 833 -114
rect 895 114 929 130
rect 895 -130 929 -114
rect 991 114 1025 130
rect 991 -130 1025 -114
rect 1087 114 1121 130
rect 1087 -130 1121 -114
rect 1183 114 1217 130
rect 1183 -130 1217 -114
rect 1279 114 1313 130
rect 1279 -130 1313 -114
rect -1281 -207 -1265 -173
rect -1231 -207 -1215 -173
rect -1089 -207 -1073 -173
rect -1039 -207 -1023 -173
rect -897 -207 -881 -173
rect -847 -207 -831 -173
rect -705 -207 -689 -173
rect -655 -207 -639 -173
rect -513 -207 -497 -173
rect -463 -207 -447 -173
rect -321 -207 -305 -173
rect -271 -207 -255 -173
rect -129 -207 -113 -173
rect -79 -207 -63 -173
rect 63 -207 79 -173
rect 113 -207 129 -173
rect 255 -207 271 -173
rect 305 -207 321 -173
rect 447 -207 463 -173
rect 497 -207 513 -173
rect 639 -207 655 -173
rect 689 -207 705 -173
rect 831 -207 847 -173
rect 881 -207 897 -173
rect 1023 -207 1039 -173
rect 1073 -207 1089 -173
rect 1215 -207 1231 -173
rect 1265 -207 1281 -173
<< viali >>
rect -1313 -114 -1279 114
rect -1217 -114 -1183 114
rect -1121 -114 -1087 114
rect -1025 -114 -991 114
rect -929 -114 -895 114
rect -833 -114 -799 114
rect -737 -114 -703 114
rect -641 -114 -607 114
rect -545 -114 -511 114
rect -449 -114 -415 114
rect -353 -114 -319 114
rect -257 -114 -223 114
rect -161 -114 -127 114
rect -65 -114 -31 114
rect 31 -114 65 114
rect 127 -114 161 114
rect 223 -114 257 114
rect 319 -114 353 114
rect 415 -114 449 114
rect 511 -114 545 114
rect 607 -114 641 114
rect 703 -114 737 114
rect 799 -114 833 114
rect 895 -114 929 114
rect 991 -114 1025 114
rect 1087 -114 1121 114
rect 1183 -114 1217 114
rect 1279 -114 1313 114
<< metal1 >>
rect -1319 114 -1273 126
rect -1319 -114 -1313 114
rect -1279 -114 -1273 114
rect -1319 -126 -1273 -114
rect -1223 114 -1177 126
rect -1223 -114 -1217 114
rect -1183 -114 -1177 114
rect -1223 -126 -1177 -114
rect -1127 114 -1081 126
rect -1127 -114 -1121 114
rect -1087 -114 -1081 114
rect -1127 -126 -1081 -114
rect -1031 114 -985 126
rect -1031 -114 -1025 114
rect -991 -114 -985 114
rect -1031 -126 -985 -114
rect -935 114 -889 126
rect -935 -114 -929 114
rect -895 -114 -889 114
rect -935 -126 -889 -114
rect -839 114 -793 126
rect -839 -114 -833 114
rect -799 -114 -793 114
rect -839 -126 -793 -114
rect -743 114 -697 126
rect -743 -114 -737 114
rect -703 -114 -697 114
rect -743 -126 -697 -114
rect -647 114 -601 126
rect -647 -114 -641 114
rect -607 -114 -601 114
rect -647 -126 -601 -114
rect -551 114 -505 126
rect -551 -114 -545 114
rect -511 -114 -505 114
rect -551 -126 -505 -114
rect -455 114 -409 126
rect -455 -114 -449 114
rect -415 -114 -409 114
rect -455 -126 -409 -114
rect -359 114 -313 126
rect -359 -114 -353 114
rect -319 -114 -313 114
rect -359 -126 -313 -114
rect -263 114 -217 126
rect -263 -114 -257 114
rect -223 -114 -217 114
rect -263 -126 -217 -114
rect -167 114 -121 126
rect -167 -114 -161 114
rect -127 -114 -121 114
rect -167 -126 -121 -114
rect -71 114 -25 126
rect -71 -114 -65 114
rect -31 -114 -25 114
rect -71 -126 -25 -114
rect 25 114 71 126
rect 25 -114 31 114
rect 65 -114 71 114
rect 25 -126 71 -114
rect 121 114 167 126
rect 121 -114 127 114
rect 161 -114 167 114
rect 121 -126 167 -114
rect 217 114 263 126
rect 217 -114 223 114
rect 257 -114 263 114
rect 217 -126 263 -114
rect 313 114 359 126
rect 313 -114 319 114
rect 353 -114 359 114
rect 313 -126 359 -114
rect 409 114 455 126
rect 409 -114 415 114
rect 449 -114 455 114
rect 409 -126 455 -114
rect 505 114 551 126
rect 505 -114 511 114
rect 545 -114 551 114
rect 505 -126 551 -114
rect 601 114 647 126
rect 601 -114 607 114
rect 641 -114 647 114
rect 601 -126 647 -114
rect 697 114 743 126
rect 697 -114 703 114
rect 737 -114 743 114
rect 697 -126 743 -114
rect 793 114 839 126
rect 793 -114 799 114
rect 833 -114 839 114
rect 793 -126 839 -114
rect 889 114 935 126
rect 889 -114 895 114
rect 929 -114 935 114
rect 889 -126 935 -114
rect 985 114 1031 126
rect 985 -114 991 114
rect 1025 -114 1031 114
rect 985 -126 1031 -114
rect 1081 114 1127 126
rect 1081 -114 1087 114
rect 1121 -114 1127 114
rect 1081 -126 1127 -114
rect 1177 114 1223 126
rect 1177 -114 1183 114
rect 1217 -114 1223 114
rect 1177 -126 1223 -114
rect 1273 114 1319 126
rect 1273 -114 1279 114
rect 1313 -114 1319 114
rect 1273 -126 1319 -114
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.26 l 0.15 m 1 nf 27 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
