* SPICE3 file created from cp1_buffer_5stage.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_HRDN5X a_n129_n130# a_n369_n42# a_543_64# a_63_n130#
+ a_159_64# a_n417_64# a_687_n42# a_303_n42# a_n561_n42# a_n321_n130# a_n749_n42#
+ a_639_n130# a_n81_n42# a_399_n42# a_n273_n42# a_15_n42# a_447_n130# a_n609_64# a_591_n42#
+ a_207_n42# a_n465_n42# a_351_64# a_255_n130# a_n33_64# a_n225_64# a_n705_n130# a_n177_n42#
+ a_n657_n42# a_495_n42# a_111_n42# a_n513_n130# VSUBS
X0 a_303_n42# a_255_n130# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_591_n42# a_543_64# a_495_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_207_n42# a_159_64# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_399_n42# a_351_64# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_495_n42# a_447_n130# a_399_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_687_n42# a_639_n130# a_591_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n561_n42# a_n609_64# a_n657_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n657_n42# a_n705_n130# a_n749_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X8 a_n465_n42# a_n513_n130# a_n561_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n369_n42# a_n417_64# a_n465_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n273_n42# a_n321_n130# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n81_n42# a_n129_n130# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n177_n42# a_n225_64# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MH6KF8 c1_n1046_n900# m3_n1086_n940# VSUBS
X0 c1_n1046_n900# m3_n1086_n940# sky130_fd_pr__cap_mim_m3_1 l=9 w=9
C0 c1_n1046_n900# m3_n1086_n940# 7.78f
C1 m3_n1086_n940# VSUBS 3.31f
.ends

.subckt nmos_dnw3 vin out1 out2 clk clkb vs VSUBS
X0 clkb clk vin vs sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.126 ps=1.44 w=0.42 l=0.15
X1 vin clkb clk vs sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.13 ps=1.46 w=0.42 l=0.15
X2 out2 clk vin vs sky130_fd_pr__nfet_01v8 ad=1.65 pd=7.1 as=0.945 ps=3.63 w=3 l=1
X3 vin clkb out1 vs sky130_fd_pr__nfet_01v8 ad=0.945 pd=3.63 as=1.65 ps=7.1 w=3 l=1
C0 vs VSUBS 6.64f
.ends

.subckt sky130_fd_pr__pfet_01v8_FBZ64Q a_n81_n126# a_399_n126# a_351_n223# a_n417_n223#
+ a_207_n126# a_n225_n223# a_n461_n126# a_n369_n126# a_63_157# a_303_n126# a_255_157#
+ a_n33_n223# a_15_n126# a_n177_n126# a_n129_157# a_111_n126# w_n497_n226# a_n273_n126#
+ a_159_n223# a_n321_157# VSUBS
X0 a_n273_n126# a_n321_157# a_n369_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_207_n126# a_159_n223# a_111_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2 a_n177_n126# a_n225_n223# a_n273_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 a_111_n126# a_63_157# a_15_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_399_n126# a_351_n223# a_303_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_n81_n126# a_n129_157# a_n177_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X6 a_15_n126# a_n33_n223# a_n81_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X7 a_n369_n126# a_n417_n223# a_n461_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X8 a_303_n126# a_255_157# a_207_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_5ACVEW a_n129_n130# a_63_n130# a_n81_n42# a_15_n42#
+ a_n173_n42# a_n33_64# a_111_n42# VSUBS
X0 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n81_n42# a_n129_n130# a_n173_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGLN5 a_n129_n130# a_n369_n42# a_1215_n130# a_543_64#
+ a_63_n130# a_159_64# a_n1089_n130# a_n849_n42# a_n417_64# a_n801_64# a_687_n42#
+ a_303_n42# a_1167_n42# a_n561_n42# a_n321_n130# a_n1041_n42# a_639_n130# a_n1185_64#
+ a_1023_n130# a_n1281_n130# a_n81_n42# a_399_n42# a_879_n42# a_n273_n42# a_735_64#
+ a_n753_n42# a_15_n42# a_n897_n130# a_n1233_n42# a_831_n130# a_447_n130# a_n609_64#
+ a_1071_n42# a_591_n42# a_1119_64# a_n993_64# a_207_n42# a_n465_n42# a_n945_n42#
+ a_351_64# a_783_n42# a_255_n130# a_n33_64# a_n225_64# a_n705_n130# a_1263_n42# a_927_64#
+ a_n177_n42# a_n657_n42# a_n1325_n42# a_n1137_n42# a_495_n42# a_111_n42# a_975_n42#
+ a_n513_n130# VSUBS
X0 a_303_n42# a_255_n130# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_591_n42# a_543_64# a_495_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_207_n42# a_159_64# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_399_n42# a_351_64# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_495_n42# a_447_n130# a_399_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_687_n42# a_639_n130# a_591_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_783_n42# a_735_64# a_687_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_975_n42# a_927_64# a_879_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n1041_n42# a_n1089_n130# a_n1137_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_879_n42# a_831_n130# a_783_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n1233_n42# a_n1281_n130# a_n1325_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X11 a_n1137_n42# a_n1185_64# a_n1233_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n561_n42# a_n609_64# a_n657_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1071_n42# a_1023_n130# a_975_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1263_n42# a_1215_n130# a_1167_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n945_n42# a_n993_64# a_n1041_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n753_n42# a_n801_64# a_n849_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n657_n42# a_n705_n130# a_n753_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n465_n42# a_n513_n130# a_n561_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n369_n42# a_n417_64# a_n465_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_1167_n42# a_1119_64# a_1071_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n849_n42# a_n897_n130# a_n945_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n273_n42# a_n321_n130# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n81_n42# a_n129_n130# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n177_n42# a_n225_64# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_VR4B8J a_1119_157# a_783_n126# a_n81_n126# a_n849_n126#
+ a_399_n126# a_n1041_n126# a_351_157# a_495_n126# a_n945_n126# a_n33_157# a_n129_n223#
+ a_n513_n223# a_1215_n223# a_63_n223# a_n1089_n223# a_n225_157# a_591_n126# a_n657_n126#
+ a_207_n126# a_543_157# a_n1325_n126# a_n369_n126# a_n753_n126# a_n321_n223# a_303_n126#
+ a_1023_n223# a_639_n223# a_n1281_n223# a_n417_157# a_n465_n126# a_1167_n126# a_735_157#
+ a_15_n126# a_n561_n126# a_n993_157# a_n177_n126# a_n897_n223# w_n1361_n226# a_1263_n126#
+ a_879_n126# a_111_n126# a_831_n223# a_n609_157# a_447_n223# a_n273_n126# a_n1137_n126#
+ a_975_n126# a_927_157# a_n1185_157# a_n1233_n126# a_n801_157# a_1071_n126# a_687_n126#
+ a_255_n223# a_n705_n223# a_159_157# VSUBS
X0 a_n273_n126# a_n321_n223# a_n369_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_n1233_n126# a_n1281_n223# a_n1325_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2 a_591_n126# a_543_157# a_495_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 a_n849_n126# a_n897_n223# a_n945_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_207_n126# a_159_157# a_111_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_n177_n126# a_n225_157# a_n273_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X6 a_n1137_n126# a_n1185_157# a_n1233_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X7 a_495_n126# a_447_n223# a_399_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X8 a_n561_n126# a_n609_157# a_n657_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X9 a_111_n126# a_63_n223# a_15_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X10 a_783_n126# a_735_157# a_687_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X11 a_1071_n126# a_1023_n223# a_975_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X12 a_399_n126# a_351_157# a_303_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X13 a_n465_n126# a_n513_n223# a_n561_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X14 a_687_n126# a_639_n223# a_591_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X15 a_n753_n126# a_n801_157# a_n849_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X16 a_975_n126# a_927_157# a_879_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X17 a_n81_n126# a_n129_n223# a_n177_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X18 a_15_n126# a_n33_157# a_n81_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X19 a_1263_n126# a_1215_n223# a_1167_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X20 a_n1041_n126# a_n1089_n223# a_n1137_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X21 a_n369_n126# a_n417_157# a_n465_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X22 a_n657_n126# a_n705_n223# a_n753_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X23 a_879_n126# a_831_n223# a_783_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X24 a_n945_n126# a_n993_157# a_n1041_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X25 a_1167_n126# a_1119_157# a_1071_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X26 a_303_n126# a_255_n223# a_207_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
C0 w_n1361_n226# VSUBS 3.67f
.ends

.subckt inverter_27x m1_n804_1398# m1_540_1398# m1_156_1398# m1_n36_1398# m1_732_1398#
+ m1_n1102_1398# m1_348_1398# m1_n1188_1398# m1_n996_1398# m1_n228_1398# m1_n1188_1912#
+ m1_924_1398# m1_1309_1398# a_n1158_1658# m1_n420_1398# m1_1116_1398# w_1358_2036#
+ m1_n612_1398# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1658# m1_n228_1398# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# a_n1158_1658# a_n1158_1658#
+ m1_n1102_1398# m1_n1102_1398# m1_1309_1398# m1_n420_1398# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_540_1398#
+ m1_n1102_1398# m1_n1102_1398# a_n1158_1658# m1_n612_1398# m1_156_1398# a_n1158_1658#
+ m1_n1102_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_732_1398#
+ a_n1158_1658# a_n1158_1658# m1_348_1398# m1_n1102_1398# m1_n804_1398# a_n1158_1658#
+ m1_924_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# m1_n36_1398# m1_n1102_1398# m1_n1188_1398# m1_n996_1398# m1_n1102_1398#
+ m1_n1102_1398# m1_1116_1398# a_n1158_1658# VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1658# m1_n1188_1912# m1_1309_1398# m1_1309_1398#
+ m1_n1188_1912# m1_1309_1398# a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ m1_n1188_1912# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ a_n1158_1658# m1_n1188_1912# a_n1158_1658# w_1358_2036# m1_1309_1398# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_1309_1398# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# a_n1158_1658# m1_1309_1398# a_n1158_1658# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
C0 a_n1158_1658# VSUBS 6.39f
C1 w_1358_2036# VSUBS 3.69f
.ends

.subckt sky130_fd_pr__nfet_01v8_KMMFCM a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_29EZRJ a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_FL984Q a_n81_n126# a_n33_157# a_n129_n223# a_63_n223#
+ a_n173_n126# a_15_n126# a_111_n126# w_n209_n226# VSUBS
X0 a_111_n126# a_63_n223# a_15_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_n81_n126# a_n129_n223# a_n173_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2 a_15_n126# a_n33_157# a_n81_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_FXZ64Q a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_D4CDWR a_n369_n42# a_n225_n130# a_303_n42# a_n81_n42#
+ a_399_n42# a_n33_n130# a_n273_n42# a_n461_n42# a_15_n42# a_n321_64# a_207_n42# a_159_n130#
+ a_n177_n42# a_351_n130# a_255_64# a_n417_n130# a_111_n42# a_n129_64# a_63_64# VSUBS
X0 a_303_n42# a_255_64# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_207_n42# a_159_n130# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_399_n42# a_351_n130# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n369_n42# a_n417_n130# a_n461_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4 a_15_n42# a_n33_n130# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_111_n42# a_63_64# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n273_n42# a_n321_64# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n81_n42# a_n129_64# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n177_n42# a_n225_n130# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_DQBD8A a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt clock clk_in vdd gnd clk clkb
Xsky130_fd_pr__pfet_01v8_FBZ64Q_0 vdd a_3246_118# a_2402_572# a_2402_572# a_3246_118#
+ a_2402_572# vdd a_3246_118# a_2402_572# vdd a_2402_572# a_2402_572# a_3246_118#
+ a_3246_118# a_2402_572# vdd vdd vdd a_2402_572# a_2402_572# gnd sky130_fd_pr__pfet_01v8_FBZ64Q
Xsky130_fd_pr__nfet_01v8_5ACVEW_0 a_344_n986# a_344_n986# a_2402_572# gnd gnd a_344_n986#
+ a_2402_572# gnd sky130_fd_pr__nfet_01v8_5ACVEW
Xinverter_27x_0 clk clk clk clk clk gnd clk clk clk clk vdd clk clk a_3246_118# clk
+ clk vdd clk gnd inverter_27x
Xsky130_fd_pr__nfet_01v8_KMMFCM_0 a_134_122# clk_in gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_1 a_416_120# a_344_102# sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42#
+ gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_2 sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42# a_134_122#
+ gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__pfet_01v8_29EZRJ_0 vdd vdd a_134_122# clk_in gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FL984Q_0 a_2402_572# a_344_n986# a_344_n986# a_344_n986#
+ vdd vdd a_2402_572# vdd gnd sky130_fd_pr__pfet_01v8_FL984Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 vdd vdd a_1230_122# m1_998_498# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_1 a_416_120# vdd vdd a_344_102# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 vdd vdd a_1430_122# a_1230_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_2 vdd vdd a_416_120# a_134_122# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_2 vdd vdd a_344_n986# a_1430_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_3 vdd vdd m1_998_498# a_786_n2# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__nfet_01v8_D4CDWR_0 a_3246_118# a_2402_572# gnd gnd a_3246_118# a_2402_572#
+ gnd gnd a_3246_118# a_2402_572# a_3246_118# a_2402_572# a_3246_118# a_2402_572#
+ a_2402_572# a_2402_572# gnd a_2402_572# a_2402_572# gnd sky130_fd_pr__nfet_01v8_D4CDWR
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 m1_998_498# a_786_n2# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 a_1230_122# m1_998_498# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_2 a_1430_122# a_1230_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_3 a_344_n986# a_1430_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
X0 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 vdd a_344_102# a_2020_n482# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X5 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X7 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X9 a_786_n912# a_586_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X10 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X11 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X12 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X13 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X17 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X20 a_286_n478# clk_in gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.15
X21 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X22 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X24 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_586_n2# a_416_120# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X27 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X28 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X30 a_786_n912# a_586_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X31 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X32 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 vdd a_344_n986# a_286_n960# vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.183 ps=1.55 w=1.26 l=0.15
X34 a_344_102# a_1394_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X35 a_992_n918# a_786_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X36 a_1192_n918# a_992_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X37 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X38 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X39 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1394_n918# a_1192_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X42 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X43 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X46 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X48 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X49 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X51 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X52 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_586_n912# a_286_n960# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X54 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X55 a_586_n2# a_416_120# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X56 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X57 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X58 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X59 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X61 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X63 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X66 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X68 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_786_n2# a_586_n2# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X72 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_286_n960# clk_in vdd vdd sky130_fd_pr__pfet_01v8 ad=0.183 pd=1.55 as=0.365 ps=3.1 w=1.26 l=0.15
X74 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X75 a_286_n960# a_344_n986# a_286_n478# gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.15
X76 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X77 a_586_n912# a_286_n960# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X78 a_1394_n918# a_1192_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X79 a_1192_n918# a_992_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X80 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X81 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X82 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X83 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X84 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X85 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X86 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X87 a_344_102# a_1394_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X88 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X89 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X90 gnd a_344_102# a_2020_n482# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X91 a_992_n918# a_786_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X92 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X93 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X94 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X95 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X96 a_786_n2# a_586_n2# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X97 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
C0 a_2432_n962# clkb 2.67f
C1 vdd a_2432_n962# 7.04f
C2 vdd clkb 7.31f
C3 vdd a_2020_n482# 2.66f
C4 clkb gnd 5.1f
C5 a_2432_n962# gnd 8.71f
C6 a_2020_n482# gnd 2.57f
C7 vdd gnd 26.1f
C8 a_344_102# gnd 2.81f
C9 a_2402_572# gnd 2.31f
C10 a_344_n986# gnd 2.43f
C11 a_3246_118# gnd 6.79f
.ends

.subckt buffer_digital m1_304_98# a_n274_130# sky130_fd_pr__pfet_01v8_FXZ64Q_1/VSUBS
+ w_n192_202#
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 w_n192_202# w_n192_202# a_116_148# a_n274_130# sky130_fd_pr__pfet_01v8_FXZ64Q_1/VSUBS
+ sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 w_n192_202# w_n192_202# m1_304_98# a_116_148# sky130_fd_pr__pfet_01v8_FXZ64Q_1/VSUBS
+ sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 a_116_148# a_n274_130# sky130_fd_pr__pfet_01v8_FXZ64Q_1/VSUBS
+ sky130_fd_pr__pfet_01v8_FXZ64Q_1/VSUBS sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 m1_304_98# a_116_148# sky130_fd_pr__pfet_01v8_FXZ64Q_1/VSUBS
+ sky130_fd_pr__pfet_01v8_FXZ64Q_1/VSUBS sky130_fd_pr__nfet_01v8_DQBD8A
.ends

.subckt sky130_fd_pr__pfet_01v8_4ZKXAA a_63_n42# a_n417_n42# a_303_n139# w_n545_n142#
+ a_255_n42# a_n465_n139# a_n129_n42# a_111_n139# a_447_n42# a_n273_n139# a_n177_73#
+ a_n321_n42# a_207_73# a_n509_n42# a_159_n42# a_15_73# a_n81_n139# a_351_n42# a_n33_n42#
+ a_n369_73# a_n225_n42# a_399_73# VSUBS
X0 a_n33_n42# a_n81_n139# a_n129_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_351_n42# a_303_n139# a_255_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n139# a_63_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_73# a_159_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_447_n42# a_399_73# a_351_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_73# a_n417_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n225_n42# a_n273_n139# a_n321_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n139# a_n509_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X8 a_n129_n42# a_n177_73# a_n225_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_63_n42# a_15_73# a_n33_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_9LGCGE a_15_n130# a_n561_n130# a_63_n42# a_n989_n42#
+ a_n177_n130# a_n417_n42# a_n465_64# a_255_n42# a_495_64# a_735_n42# a_n129_n42#
+ a_n609_n42# a_111_64# a_447_n42# a_927_n42# a_783_n130# a_n321_n42# a_399_n130#
+ a_n657_64# a_n801_n42# a_687_64# a_n945_n130# a_159_n42# a_639_n42# a_n513_n42#
+ a_n897_n42# a_591_n130# a_n81_64# a_n273_64# a_351_n42# a_207_n130# a_303_64# a_n33_n42#
+ a_831_n42# a_n369_n130# a_n753_n130# a_n849_64# a_n225_n42# a_n705_n42# a_879_64#
+ a_543_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n897_n42# a_n945_n130# a_n989_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_49FP49 a_63_n42# a_n989_n42# a_n369_n139# a_n753_n139#
+ a_n417_n42# a_687_73# w_n1025_n142# a_255_n42# a_735_n42# a_n81_73# a_n273_73# a_n129_n42#
+ a_15_n139# a_n561_n139# a_303_73# a_n609_n42# a_n177_n139# a_n849_73# a_447_n42#
+ a_927_n42# a_n321_n42# a_879_73# a_n801_n42# a_159_n42# a_639_n42# a_n465_73# a_n513_n42#
+ a_n897_n42# a_783_n139# a_495_73# a_399_n139# a_351_n42# a_n33_n42# a_831_n42# a_n945_n139#
+ a_n225_n42# a_n705_n42# a_111_73# a_591_n139# a_543_n42# a_207_n139# a_n657_73#
+ VSUBS
X0 a_927_n42# a_879_73# a_831_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_73# a_n129_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_73# a_255_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_73# a_63_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n139# a_159_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_n139# a_351_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_543_n42# a_495_73# a_447_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_639_n42# a_591_n139# a_543_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_73# a_639_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n139# a_735_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n801_n42# a_n849_73# a_n897_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n513_n42# a_n561_n139# a_n609_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n321_n42# a_n369_n139# a_n417_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n225_n42# a_n273_73# a_n321_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n897_n42# a_n945_n139# a_n989_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X15 a_n705_n42# a_n753_n139# a_n801_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n609_n42# a_n657_73# a_n705_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n417_n42# a_n465_73# a_n513_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n139# a_n225_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_63_n42# a_15_n139# a_n33_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC45 a_63_n42# a_15_64# a_n417_n42# a_111_n130#
+ a_n273_n130# a_255_n42# a_n129_n42# a_n369_64# a_399_64# a_447_n42# a_n81_n130#
+ a_n321_n42# a_n509_n42# a_159_n42# a_351_n42# a_n33_n42# a_303_n130# a_n225_n42#
+ a_n177_64# a_207_64# a_n465_n130# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_n130# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_64# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n321_n42# a_n369_64# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n130# a_n509_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X8 a_n225_n42# a_n273_n130# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt buffer m1_n1188_2032# a_1504_1398# m1_n1188_1271# m5_n1320_776# a_n1158_1778#
+ a_1504_1860# a_1596_1398# w_1358_2156# m4_n1330_2222# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1778# m1_n1188_1271# a_n1158_1778# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778#
+ a_1436_1552# a_1436_1552# m1_n1188_1271# m1_n1188_1271# a_n1158_1778# a_1436_1552#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# m1_n1188_1271#
+ a_1436_1552# a_1436_1552# a_n1158_1778# m1_n1188_1271# m1_n1188_1271# a_n1158_1778#
+ a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# m1_n1188_1271#
+ a_n1158_1778# a_n1158_1778# m1_n1188_1271# a_1436_1552# m1_n1188_1271# a_n1158_1778#
+ m1_n1188_1271# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552#
+ a_n1158_1778# m1_n1188_1271# a_1436_1552# m1_n1188_1271# m1_n1188_1271# a_1436_1552#
+ a_1436_1552# m1_n1188_1271# a_n1158_1778# VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1778# m1_n1188_2032# a_1436_1552# a_1436_1552#
+ m1_n1188_2032# a_1436_1552# a_n1158_1778# a_1436_1552# m1_n1188_2032# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ m1_n1188_2032# a_1436_1552# m1_n1188_2032# a_n1158_1778# m1_n1188_2032# m1_n1188_2032#
+ m1_n1188_2032# a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ a_n1158_1778# a_1436_1552# m1_n1188_2032# a_n1158_1778# m1_n1188_2032# m1_n1188_2032#
+ a_n1158_1778# m1_n1188_2032# a_n1158_1778# w_1358_2156# a_1436_1552# a_1436_1552#
+ a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# m1_n1188_2032#
+ m1_n1188_2032# a_n1158_1778# a_n1158_1778# a_1436_1552# a_n1158_1778# a_1436_1552#
+ a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
X0 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X6 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X8 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X11 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X12 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X15 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X16 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X17 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X20 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X21 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X24 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X27 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X30 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X32 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X35 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X36 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X38 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X39 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X43 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X45 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X46 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X48 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X49 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X50 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X53 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
C0 a_1504_1860# a_1596_1398# 6.79f
C1 a_1436_1552# w_1358_2156# 2.61f
C2 a_1596_1398# a_1504_1398# 2.65f
C3 a_1436_1552# a_1596_1398# 2.21f
C4 m5_n1320_776# VSUBS 2.52f
C5 a_n1158_1778# VSUBS 7.08f
C6 a_1436_1552# VSUBS 8.93f
C7 w_1358_2156# VSUBS 5.14f
.ends

.subckt sky130_fd_pr__pfet_01v8_X4L24Q a_n33_n126# w_n353_n226# a_n317_n126# a_n177_157#
+ a_159_n126# a_111_n223# a_n273_n223# a_255_n126# a_n129_n126# a_n81_n223# a_63_n126#
+ a_n225_n126# a_15_157# a_207_157# VSUBS
X0 a_159_n126# a_111_n223# a_63_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_n225_n126# a_n273_n223# a_n317_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2 a_63_n126# a_15_157# a_n33_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 a_n129_n126# a_n177_157# a_n225_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_n33_n126# a_n81_n223# a_n129_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_255_n126# a_207_157# a_159_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_XJUN3E a_63_n42# a_15_64# a_111_n130# a_n273_n130#
+ a_255_n42# a_n129_n42# a_n317_n42# a_n81_n130# a_159_n42# a_n33_n42# a_n225_n42#
+ a_n177_64# a_207_64# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n225_n42# a_n273_n130# a_n317_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt and_gate a_514_134# w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206#
+ m1_748_n50#
Xsky130_fd_pr__pfet_01v8_X4L24Q_0 w_n260_286# w_n260_286# m1_748_n50# a_n78_396# w_n260_286#
+ a_n78_396# a_n78_396# m1_748_n50# m1_748_n50# a_n78_396# m1_748_n50# w_n260_286#
+ a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q
Xsky130_fd_pr__nfet_01v8_XJUN3E_0 m1_748_n50# a_n78_396# a_n78_396# a_n78_396# m1_748_n50#
+ m1_748_n50# m1_748_n50# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__nfet_01v8_XJUN3E
X0 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.57 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_n78_396# a_514_134# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X6 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 w_n260_286# a_514_134# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.195 ps=1.57 w=1.26 l=0.15
X8 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X9 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X10 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X11 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 a_n78_396# w_n260_286# 3.02f
C1 a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 2.46f
C2 w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 6.96f
.ends

.subckt buffer_and_gate in1 clk out gnd vdd
Xbuffer_0 vdd gnd gnd gnd clk vdd m1_5444_838# vdd vdd gnd buffer
Xand_gate_0 m1_5444_838# vdd gnd in1 out and_gate
C0 in1 0 2.5f
C1 and_gate_0/a_n78_396# 0 2.34f
C2 clk 0 7.7f
C3 buffer_0/a_1436_1552# 0 8.93f
C4 vdd 0 17.7f
C5 gnd 0 7.18f
.ends

.subckt capacito7 a_2858_n174# sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142# a_5270_n124#
+ m3_7758_166# buffer_and_gate_0/clk sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142#
+ m1_6370_n278# buffer_and_gate_0/gnd buffer_and_gate_0/vdd m1_602_n334# m2_n739_1036#
Xbuffer_digital_0 buffer_and_gate_0/in1 m2_n739_1036# buffer_and_gate_0/gnd buffer_and_gate_0/vdd
+ buffer_digital
Xsky130_fd_pr__pfet_01v8_4ZKXAA_0 m1_6370_n278# m1_6370_n278# buffer_and_gate_0/gnd
+ sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142# m1_6370_n278# buffer_and_gate_0/gnd
+ m1_6370_n278# buffer_and_gate_0/gnd m1_6370_n278# buffer_and_gate_0/gnd buffer_and_gate_0/gnd
+ m1_6370_n278# buffer_and_gate_0/gnd m1_6370_n278# m1_6370_n278# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd m1_6370_n278# m1_6370_n278# buffer_and_gate_0/gnd m1_6370_n278#
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__nfet_01v8_9LGCGE_0 a_2858_n174# a_2858_n174# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd a_2858_n174# buffer_and_gate_0/gnd a_2858_n174# buffer_and_gate_0/gnd
+ a_2858_n174# buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_2858_n174#
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_2858_n174# buffer_and_gate_0/gnd a_2858_n174#
+ a_2858_n174# buffer_and_gate_0/gnd a_2858_n174# a_2858_n174# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_2858_n174# a_2858_n174#
+ a_2858_n174# buffer_and_gate_0/gnd a_2858_n174# a_2858_n174# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd a_2858_n174# a_2858_n174# a_2858_n174# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd a_2858_n174# buffer_and_gate_0/gnd buffer_and_gate_0/gnd sky130_fd_pr__nfet_01v8_9LGCGE
Xsky130_fd_pr__pfet_01v8_49FP49_0 m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd m1_602_n334# buffer_and_gate_0/gnd sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142#
+ m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd buffer_and_gate_0/gnd m1_602_n334#
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd m1_602_n334# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd m1_602_n334# m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd
+ m1_602_n334# m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd m1_602_n334# m1_602_n334#
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd m1_602_n334# m1_602_n334#
+ m1_602_n334# buffer_and_gate_0/gnd m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd m1_602_n334# buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd
+ sky130_fd_pr__pfet_01v8_49FP49
Xsky130_fd_pr__nfet_01v8_NJGC45_0 buffer_and_gate_0/gnd a_5270_n124# buffer_and_gate_0/gnd
+ a_5270_n124# a_5270_n124# buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_5270_n124#
+ a_5270_n124# buffer_and_gate_0/gnd a_5270_n124# buffer_and_gate_0/gnd buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_5270_n124# buffer_and_gate_0/gnd
+ a_5270_n124# a_5270_n124# a_5270_n124# buffer_and_gate_0/gnd sky130_fd_pr__nfet_01v8_NJGC45
Xbuffer_and_gate_0 buffer_and_gate_0/in1 buffer_and_gate_0/clk buffer_and_gate_0/out
+ buffer_and_gate_0/gnd buffer_and_gate_0/vdd buffer_and_gate
X0 buffer_and_gate_0/out m3_7758_166# sky130_fd_pr__cap_mim_m3_1 l=7.99 w=7.97
C0 a_2858_n174# buffer_and_gate_0/gnd 2.03f
C1 buffer_and_gate_0/in1 m2_n739_1036# 2.94f
C2 m3_7758_166# 0 2.32f
C3 buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C4 buffer_and_gate_0/clk 0 7.7f
C5 buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C6 buffer_and_gate_0/vdd 0 18.4f
C7 buffer_and_gate_0/gnd 0 8.14f
C8 a_5270_n124# 0 2.36f
C9 a_2858_n174# 0 4.67f
C10 buffer_and_gate_0/in1 0 2.66f
.ends

.subckt capacitor_8 capacitor_7_0/a_5270_n124# capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/vdd
+ capacitor_7_0/buffer_and_gate_0/clk capacitor_7_0/a_2858_n174# w_7118_n356# w_1380_n364#
+ VSUBS capacitor_7_0/m2_n739_1036#
Xcapacitor_7_0 capacitor_7_0/a_2858_n174# w_7118_n356# capacitor_7_0/a_5270_n124#
+ capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/clk w_1380_n364# w_7118_n356#
+ VSUBS capacitor_7_0/buffer_and_gate_0/vdd w_1380_n364# capacitor_7_0/m2_n739_1036#
+ capacito7
C0 capacitor_7_0/m3_7758_166# 0 2.32f
C1 capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C2 capacitor_7_0/buffer_and_gate_0/clk 0 7.7f
C3 capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C4 capacitor_7_0/buffer_and_gate_0/vdd 0 18.5f
C5 VSUBS 0 7.98f
C6 capacitor_7_0/a_5270_n124# 0 2.36f
C7 w_1380_n364# 0 3.28f
C8 capacitor_7_0/a_2858_n174# 0 4.67f
C9 capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
.ends

.subckt capacitors_1 clk1 in1 capacitor_8_0/capacitor_7_0/a_2858_n174# capacitor_8_0/capacitor_7_0/a_5270_n124#
+ capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk capacitor_8_0/capacitor_7_0/buffer_and_gate_0/vdd
+ m1_7096_n308# capacitor_8_0/w_1380_n364# VSUBS
Xcapacitor_8_0 capacitor_8_0/capacitor_7_0/a_5270_n124# clk1 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/vdd
+ capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk capacitor_8_0/capacitor_7_0/a_2858_n174#
+ m1_7096_n308# capacitor_8_0/w_1380_n364# VSUBS in1 capacitor_8
C0 VSUBS capacitor_8_0/capacitor_7_0/buffer_and_gate_0/vdd 2.84f
C1 clk1 0 2.38f
C2 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C3 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk 0 8.49f
C4 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C5 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/vdd 0 18.5f
C6 VSUBS 0 7.98f
C7 capacitor_8_0/capacitor_7_0/a_5270_n124# 0 2.36f
C8 capacitor_8_0/w_1380_n364# 0 3.28f
C9 capacitor_8_0/capacitor_7_0/a_2858_n174# 0 4.67f
C10 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
.ends

.subckt sky130_fd_pr__pfet_01v8_4RPJ49 a_2031_73# a_1887_n42# a_3615_n42# a_3183_73#
+ a_n3729_73# a_n2529_n42# a_1503_n42# a_63_n42# a_n753_n139# a_n3393_n42# a_n369_n139#
+ a_n1425_73# a_n1281_n42# a_n2961_73# a_687_73# a_n2577_73# a_n417_n42# a_2367_n42#
+ a_n1761_n42# a_n3009_n42# a_n2673_n139# a_2847_n42# a_n2289_n139# a_n3633_n139#
+ a_2607_73# a_n3249_n139# a_n1713_n139# a_3759_73# a_n1329_n139# a_255_n42# a_1455_73#
+ a_n2241_n42# a_2991_73# a_3471_n139# a_735_n42# a_1551_n139# a_3087_n139# a_1599_n42#
+ a_3327_n42# a_1167_n139# a_n2721_n42# a_n81_73# a_2511_n139# a_1215_n42# a_n273_73#
+ a_2127_n139# a_n993_n42# a_3807_n42# a_15_n139# a_303_73# a_n3585_n42# a_n129_n42#
+ a_2079_n42# a_n561_n139# a_n3345_73# a_n3201_n42# a_n1473_n42# a_n177_n139# a_n1041_73#
+ a_n609_n42# a_2559_n42# a_n2193_73# a_n1953_n42# a_n849_73# w_n3905_n142# a_n2481_n139#
+ a_n2097_n139# a_n3441_n139# a_1791_n42# a_n1521_n139# a_n3057_n139# a_2223_73# a_447_n42#
+ a_3039_n42# a_n1137_n139# a_3375_73# a_n2433_n42# a_927_n42# a_1071_73# a_n1617_73#
+ a_n2913_n42# a_3519_n42# a_975_n139# a_879_73# a_n2769_73# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n1185_n42# a_n801_n42# a_n3777_n42# a_2751_n42# a_n1665_n42#
+ a_1647_73# a_2799_73# a_3231_n42# a_159_n42# a_n2145_n42# a_n465_73# a_1983_n42#
+ a_3711_n42# a_639_n42# a_n2625_n42# a_1119_n42# a_n3537_73# a_n897_n42# a_n513_n42#
+ a_n1233_73# a_n3489_n42# a_2463_n42# a_783_n139# a_495_73# a_399_n139# a_n2385_73#
+ a_2895_n139# a_n3105_n42# a_n1377_n42# a_2943_n42# a_1935_n139# a_n1857_n42# a_351_n42#
+ a_2415_73# a_n33_n42# a_3567_73# a_831_n42# a_1695_n42# a_3423_n42# a_1263_73# a_n945_n139#
+ a_n2337_n42# a_1311_n42# a_n1809_73# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2175_n42#
+ a_n2865_n139# a_n1089_n42# a_n3825_n139# a_111_73# a_n2001_73# a_n3869_n42# a_n705_n42#
+ a_2655_n42# a_n1905_n139# a_n3153_73# a_591_n139# a_1839_73# a_n1569_n42# a_3663_n139#
+ a_1743_n139# a_3279_n139# a_543_n42# a_207_n139# a_n657_73# a_1359_n139# a_2703_n139#
+ a_3135_n42# VSUBS a_2319_n139# a_n2049_n42# a_1023_n42#
X0 a_n2241_n42# a_n2289_n139# a_n2337_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n2913_n42# a_n2961_73# a_n3009_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n2721_n42# a_n2769_73# a_n2817_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n2625_n42# a_n2673_n139# a_n2721_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n2433_n42# a_n2481_n139# a_n2529_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n2337_n42# a_n2385_73# a_n2433_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n2145_n42# a_n2193_73# a_n2241_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n2049_n42# a_n2097_n139# a_n2145_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n2817_n42# a_n2865_n139# a_n2913_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n2529_n42# a_n2577_73# a_n2625_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_2079_n42# a_2031_73# a_1983_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_2175_n42# a_2127_n139# a_2079_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_2271_n42# a_2223_73# a_2175_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_2367_n42# a_2319_n139# a_2271_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_2463_n42# a_2415_73# a_2367_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_2655_n42# a_2607_73# a_2559_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_2751_n42# a_2703_n139# a_2655_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_2943_n42# a_2895_n139# a_2847_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_2559_n42# a_2511_n139# a_2463_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_2847_n42# a_2799_73# a_2751_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_927_n42# a_879_73# a_831_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_1023_n42# a_975_n139# a_927_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n1953_n42# a_n2001_73# a_n2049_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_n1761_n42# a_n1809_73# a_n1857_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n1665_n42# a_n1713_n139# a_n1761_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n1857_n42# a_n1905_n139# a_n1953_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n1569_n42# a_n1617_73# a_n1665_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_1119_n42# a_1071_73# a_1023_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1215_n42# a_1167_n139# a_1119_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1311_n42# a_1263_73# a_1215_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_1407_n42# a_1359_n139# a_1311_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1503_n42# a_1455_73# a_1407_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_1695_n42# a_1647_73# a_1599_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1791_n42# a_1743_n139# a_1695_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1599_n42# a_1551_n139# a_1503_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_1887_n42# a_1839_73# a_1791_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_1983_n42# a_1935_n139# a_1887_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n33_n42# a_n81_73# a_n129_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_351_n42# a_303_73# a_255_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_159_n42# a_111_73# a_63_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_255_n42# a_207_n139# a_159_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_447_n42# a_399_n139# a_351_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_543_n42# a_495_73# a_447_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_639_n42# a_591_n139# a_543_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_735_n42# a_687_73# a_639_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_831_n42# a_783_n139# a_735_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_n1473_n42# a_n1521_n139# a_n1569_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_n1377_n42# a_n1425_73# a_n1473_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_n1281_n42# a_n1329_n139# a_n1377_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_n1185_n42# a_n1233_73# a_n1281_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n1089_n42# a_n1137_n139# a_n1185_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_n993_n42# a_n1041_73# a_n1089_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_n801_n42# a_n849_73# a_n897_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_n513_n42# a_n561_n139# a_n609_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_n321_n42# a_n369_n139# a_n417_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_n225_n42# a_n273_73# a_n321_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_n897_n42# a_n945_n139# a_n993_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_n705_n42# a_n753_n139# a_n801_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_n609_n42# a_n657_73# a_n705_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n417_n42# a_n465_73# a_n513_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n129_n42# a_n177_n139# a_n225_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_3327_n42# a_3279_n139# a_3231_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_3423_n42# a_3375_73# a_3327_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_3615_n42# a_3567_73# a_3519_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_3711_n42# a_3663_n139# a_3615_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_3519_n42# a_3471_n139# a_3423_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_3807_n42# a_3759_73# a_3711_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n3201_n42# a_n3249_n139# a_n3297_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_63_n42# a_15_n139# a_n33_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n3681_n42# a_n3729_73# a_n3777_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n3585_n42# a_n3633_n139# a_n3681_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n3393_n42# a_n3441_n139# a_n3489_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n3297_n42# a_n3345_73# a_n3393_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n3105_n42# a_n3153_73# a_n3201_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_n3009_n42# a_n3057_n139# a_n3105_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3231_n42# a_3183_73# a_3135_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_n3777_n42# a_n3825_n139# a_n3869_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X77 a_n3489_n42# a_n3537_73# a_n3585_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3039_n42# a_2991_73# a_2943_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3135_n42# a_3087_n139# a_3039_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 w_n3905_n142# VSUBS 6.63f
.ends

.subckt sky130_fd_pr__pfet_01v8_E9H44Q a_15_n42# a_n15_n68# w_n109_n104# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# w_n109_n104# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_9AYYDL a_n158_n300# w_n194_n362# a_100_n300# a_n100_n326#
+ VSUBS
X0 a_100_n300# a_n100_n326# a_n158_n300# w_n194_n362# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt pmos_cp1 a_168_22# m1_532_58# w_n14_n142# a_424_18# m1_14_56# VSUBS
Xsky130_fd_pr__pfet_01v8_E9H44Q_0 w_n14_n142# a_168_22# w_n14_n142# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_E9H44Q_1 a_168_22# a_424_18# w_n14_n142# w_n14_n142# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_9AYYDL_0 m1_14_56# w_n14_n142# w_n14_n142# a_168_22# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
Xsky130_fd_pr__pfet_01v8_9AYYDL_1 w_n14_n142# w_n14_n142# m1_532_58# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
C0 w_n14_n142# VSUBS 2.47f
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC8F a_15_n130# a_1887_n42# a_3615_n42# a_1647_64#
+ a_n561_n130# a_n2529_n42# a_1503_n42# a_2799_64# a_63_n42# a_n177_n130# a_n3393_n42#
+ a_n1281_n42# a_n465_64# a_n417_n42# a_2367_n42# a_n1761_n42# a_n2481_n130# a_n3009_n42#
+ a_n2097_n130# a_n3441_n130# a_2847_n42# a_n1521_n130# a_n3057_n130# a_n3537_64#
+ a_n1137_n130# a_255_n42# a_n1233_64# a_495_64# a_n2241_n42# a_n2385_64# a_975_n130#
+ a_735_n42# a_1599_n42# a_3327_n42# a_n2721_n42# a_1215_n42# a_2415_64# a_n993_n42#
+ a_3807_n42# a_3567_64# a_n3585_n42# a_n129_n42# a_2079_n42# a_1263_64# a_n3201_n42#
+ a_n1473_n42# a_n1809_64# a_n609_n42# a_2559_n42# a_n1953_n42# a_111_64# a_n2001_64#
+ a_1791_n42# a_447_n42# a_n3153_64# a_3039_n42# a_n2433_n42# a_1839_64# a_927_n42#
+ a_n2913_n42# a_3519_n42# a_783_n130# a_399_n130# a_2895_n130# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n657_64# a_n1185_n42# a_1935_n130# a_n801_n42# a_2031_64#
+ a_n3777_n42# a_2751_n42# a_3183_64# a_n1665_n42# a_n3729_64# a_n1425_64# a_687_64#
+ a_n2961_64# a_n945_n130# a_n2577_64# a_3231_n42# a_159_n42# a_n2145_n42# a_1983_n42#
+ a_3711_n42# a_2607_64# a_639_n42# a_n2625_n42# a_3759_64# a_n2865_n130# a_1119_n42#
+ a_n3825_n130# a_1455_64# a_n1905_n130# a_2991_64# a_n897_n42# a_591_n130# a_n513_n42#
+ a_n3489_n42# a_2463_n42# a_n3105_n42# a_n1377_n42# a_n81_64# a_n273_64# a_3663_n130#
+ a_3279_n130# a_2943_n42# a_1743_n130# a_207_n130# a_2703_n130# a_1359_n130# a_n1857_n42#
+ a_2319_n130# a_351_n42# a_303_64# a_n3345_64# a_n33_n42# a_831_n42# a_n1041_64#
+ a_1695_n42# a_3423_n42# a_n753_n130# a_n369_n130# a_n2193_64# a_n2337_n42# a_1311_n42#
+ a_n849_64# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2223_64# a_n2673_n130# a_2175_n42#
+ a_3375_64# a_n2289_n130# a_n3633_n130# a_n1089_n42# a_n3249_n130# a_n1713_n130#
+ a_n3869_n42# a_n705_n42# a_2655_n42# a_1071_64# a_n1329_n130# a_n1617_64# a_n1569_n42#
+ a_879_64# a_n2769_64# a_3471_n130# a_3087_n130# a_1551_n130# a_2511_n130# a_543_n42#
+ a_1167_n130# a_3135_n42# a_2127_n130# VSUBS a_n2049_n42# a_1023_n42#
X0 a_n3201_n42# a_n3249_n130# a_n3297_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n3681_n42# a_n3729_64# a_n3777_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n3585_n42# a_n3633_n130# a_n3681_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n3393_n42# a_n3441_n130# a_n3489_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n3297_n42# a_n3345_64# a_n3393_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n3105_n42# a_n3153_64# a_n3201_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n3009_n42# a_n3057_n130# a_n3105_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n3777_n42# a_n3825_n130# a_n3869_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X9 a_n3489_n42# a_n3537_64# a_n3585_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_3135_n42# a_3087_n130# a_3039_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_3231_n42# a_3183_64# a_3135_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_3039_n42# a_2991_64# a_2943_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n2241_n42# a_n2289_n130# a_n2337_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n2913_n42# a_n2961_64# a_n3009_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n2721_n42# a_n2769_64# a_n2817_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n2625_n42# a_n2673_n130# a_n2721_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n2433_n42# a_n2481_n130# a_n2529_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n2337_n42# a_n2385_64# a_n2433_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n2145_n42# a_n2193_64# a_n2241_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_n2049_n42# a_n2097_n130# a_n2145_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n2817_n42# a_n2865_n130# a_n2913_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n2529_n42# a_n2577_64# a_n2625_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2175_n42# a_2127_n130# a_2079_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_2271_n42# a_2223_64# a_2175_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2463_n42# a_2415_64# a_2367_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_2751_n42# a_2703_n130# a_2655_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_2079_n42# a_2031_64# a_1983_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_2367_n42# a_2319_n130# a_2271_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2559_n42# a_2511_n130# a_2463_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_2655_n42# a_2607_64# a_2559_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_2847_n42# a_2799_64# a_2751_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_2943_n42# a_2895_n130# a_2847_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1023_n42# a_975_n130# a_927_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_n1953_n42# a_n2001_64# a_n2049_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_n1761_n42# a_n1809_64# a_n1857_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n1665_n42# a_n1713_n130# a_n1761_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_n1857_n42# a_n1905_n130# a_n1953_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_n1569_n42# a_n1617_64# a_n1665_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1215_n42# a_1167_n130# a_1119_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1311_n42# a_1263_64# a_1215_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1503_n42# a_1455_64# a_1407_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_1791_n42# a_1743_n130# a_1695_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1119_n42# a_1071_64# a_1023_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_1407_n42# a_1359_n130# a_1311_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_1599_n42# a_1551_n130# a_1503_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1695_n42# a_1647_64# a_1599_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_1887_n42# a_1839_64# a_1791_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_1983_n42# a_1935_n130# a_1887_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n1473_n42# a_n1521_n130# a_n1569_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n1281_n42# a_n1329_n130# a_n1377_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_n1185_n42# a_n1233_64# a_n1281_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_n993_n42# a_n1041_64# a_n1089_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_n1377_n42# a_n1425_64# a_n1473_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_n1089_n42# a_n1137_n130# a_n1185_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n897_n42# a_n945_n130# a_n993_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_3327_n42# a_3279_n130# a_3231_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3423_n42# a_3375_64# a_3327_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_3615_n42# a_3567_64# a_3519_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X77 a_3711_n42# a_3663_n130# a_3615_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3519_n42# a_3471_n130# a_3423_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3807_n42# a_3759_64# a_3711_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt charge_pump1 clk_in input1 input2 in1 in5 in6 in8 g1 g2 clk clkb m1_12464_n576#
+ a_3340_18086# in4 in3 vin vdd in7 in2 gnd
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 g1 clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 g2 clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 vin input1 input2 g1 g2 vin gnd nmos_dnw3
Xclock_0 clk_in vdd gnd clk clkb clock
Xcapacitor_8_0 vdd input1 vdd clk vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 vdd clkb vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 in1 vdd vdd clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_1 input2 in1 vdd vdd clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_2 input1 in2 vdd vdd clk vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 in3 vdd vdd clk vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_4 input2 in2 vdd vdd clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_5 input2 in3 vdd vdd clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_6 input1 in4 vdd vdd clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_7 input1 in5 vdd vdd clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_8 input1 in6 vdd vdd clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_9 input1 in7 vdd vdd clk vdd vdd vdd gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 in7 vdd vdd clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_11 input2 in6 vdd vdd clkb vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 in4 vdd vdd clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_12 input2 in5 vdd vdd clkb vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clkb input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clk input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 vdd input1 26.8f
C1 vdd input2 26.5f
C2 vin clk 2.19f
C3 clk m1_12464_n576# 2.31f
C4 input2 input1 3.06f
C5 clkb m1_12464_n576# 2.21f
C6 gnd clk 2.59f
C7 vin vdd 9.14f
C8 gnd vdd 0.171p
C9 gnd input1 8.5f
C10 gnd input2 8.88f
C11 vdd clk 32.2f
C12 vdd clkb 26.2f
C13 input1 0 22.5f
C14 input2 0 22.2f
C15 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C16 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C17 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C18 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C19 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C20 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C21 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C22 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C23 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C24 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C25 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C26 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C27 m1_4341_n519# 0 3.77f
C28 m1_12659_300# 0 2.54f
C29 m1_12464_n576# 0 4.25f
C30 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C31 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C32 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C33 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C34 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C35 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C36 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C37 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C38 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C39 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C40 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C41 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C42 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C43 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C44 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C45 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C46 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C47 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C48 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C49 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C50 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C51 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C52 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C53 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C54 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C55 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C56 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C57 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C58 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C59 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C60 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C61 clkb 0 85.9f
C62 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C63 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C64 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C65 clk 0 85.1f
C66 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C67 vdd 0 0.461p
C68 gnd 0 45.3f
C69 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C70 clock_0/a_2432_n962# 0 8.68f **FLOATING
C71 clock_0/a_2020_n482# 0 2.57f **FLOATING
C72 clock_0/a_344_102# 0 2.81f
C73 clock_0/a_2402_572# 0 2.17f
C74 clock_0/a_344_n986# 0 2.38f
C75 clock_0/a_3246_118# 0 6.83f
C76 g2 0 2.34f
C77 vin 0 10.4f
.ends

.subckt sky130_fd_pr__nfet_01v8_TKGCLY a_n1425_n130# a_1887_n42# a_1503_n42# a_63_n42#
+ a_15_64# a_2127_64# a_n1281_n42# a_111_n130# a_879_n130# a_1263_n130# a_n417_n42#
+ a_2367_n42# a_2223_n130# a_n1761_n42# a_n1905_64# a_n273_n130# a_255_n42# a_n2241_n42#
+ a_735_n42# a_1599_n42# a_1935_64# a_n2429_n42# a_1215_n42# a_n2193_n130# a_n993_n42#
+ a_n1233_n130# a_n753_64# a_n369_64# a_n129_n42# a_2079_n42# a_n1473_n42# a_n609_n42#
+ a_687_n130# a_1071_n130# a_n1953_n42# a_2031_n130# a_n1521_64# a_n1137_64# a_783_64#
+ a_399_64# a_1839_n130# a_n2289_64# a_1791_n42# a_447_n42# a_927_n42# a_n81_n130#
+ a_2319_64# a_n849_n130# a_n321_n42# a_1407_n42# a_1551_64# a_2271_n42# a_1167_64#
+ a_n1185_n42# a_n801_n42# a_n1041_n130# a_n2001_n130# a_n1665_n42# a_n1809_n130#
+ a_495_n130# a_159_n42# a_n2145_n42# a_1647_n130# a_1983_n42# a_639_n42# a_n945_64#
+ a_1119_n42# a_n897_n42# a_n657_n130# a_n513_n42# a_n1377_n42# a_n1713_64# a_n1329_64#
+ a_975_64# a_n1857_n42# a_351_n42# a_n33_n42# a_n1617_n130# a_831_n42# a_1695_n42#
+ a_n2337_n42# a_1311_n42# a_303_n130# a_1743_64# a_1359_64# a_1455_n130# a_n225_n42#
+ a_2175_n42# a_n561_64# a_n1089_n42# a_n177_64# a_n705_n42# a_n465_n130# a_n1569_n42#
+ a_207_64# a_543_n42# a_591_64# a_n2097_64# a_n2385_n130# VSUBS a_n2049_n42# a_1023_n42#
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n2241_n42# a_n2289_64# a_n2337_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n2337_n42# a_n2385_n130# a_n2429_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3 a_n2145_n42# a_n2193_n130# a_n2241_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n2049_n42# a_n2097_64# a_n2145_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_2175_n42# a_2127_64# a_2079_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_2271_n42# a_2223_n130# a_2175_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_2079_n42# a_2031_n130# a_1983_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_2367_n42# a_2319_64# a_2271_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_927_n42# a_879_n130# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_1023_n42# a_975_64# a_927_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n1953_n42# a_n2001_n130# a_n2049_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n1761_n42# a_n1809_n130# a_n1857_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n1665_n42# a_n1713_64# a_n1761_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n1857_n42# a_n1905_64# a_n1953_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n1569_n42# a_n1617_n130# a_n1665_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_1215_n42# a_1167_64# a_1119_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_1311_n42# a_1263_n130# a_1215_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_1503_n42# a_1455_n130# a_1407_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_1791_n42# a_1743_64# a_1695_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_1119_n42# a_1071_n130# a_1023_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_1407_n42# a_1359_64# a_1311_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1599_n42# a_1551_64# a_1503_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_1695_n42# a_1647_n130# a_1599_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_1887_n42# a_1839_n130# a_1791_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_1983_n42# a_1935_64# a_1887_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_351_n42# a_303_n130# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_447_n42# a_399_64# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_543_n42# a_495_n130# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_735_n42# a_687_n130# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_831_n42# a_783_64# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_639_n42# a_591_64# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_n1473_n42# a_n1521_64# a_n1569_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_n1281_n42# a_n1329_64# a_n1377_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n1185_n42# a_n1233_n130# a_n1281_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_n993_n42# a_n1041_n130# a_n1089_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_n1377_n42# a_n1425_n130# a_n1473_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_n1089_n42# a_n1137_64# a_n1185_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_n321_n42# a_n369_64# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_n801_n42# a_n849_n130# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_n705_n42# a_n753_64# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_n609_n42# a_n657_n130# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_n513_n42# a_n561_64# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_n417_n42# a_n465_n130# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_n225_n42# a_n273_n130# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_n897_n42# a_n945_64# a_n993_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt nmos_decap_10 a_n2_210# m1_n10_n42# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGC45_0 m1_n10_n42# a_n2_210# m1_n10_n42# a_n2_210# a_n2_210#
+ m1_n10_n42# m1_n10_n42# a_n2_210# a_n2_210# m1_n10_n42# a_n2_210# m1_n10_n42# m1_n10_n42#
+ m1_n10_n42# m1_n10_n42# m1_n10_n42# a_n2_210# m1_n10_n42# a_n2_210# a_n2_210# a_n2_210#
+ VSUBS sky130_fd_pr__nfet_01v8_NJGC45
C0 a_n2_210# VSUBS 2.33f
.ends

.subckt pmos_decap_10 a_12_230# w_6_4# VSUBS
Xsky130_fd_pr__pfet_01v8_4ZKXAA_0 w_6_4# w_6_4# a_12_230# w_6_4# w_6_4# a_12_230#
+ w_6_4# a_12_230# w_6_4# a_12_230# a_12_230# w_6_4# a_12_230# w_6_4# w_6_4# a_12_230#
+ a_12_230# w_6_4# w_6_4# a_12_230# w_6_4# a_12_230# VSUBS sky130_fd_pr__pfet_01v8_4ZKXAA
.ends

.subckt cp1_buffer1 charge_pump1_0/clk_in charge_pump1_0/in3 charge_pump1_0/in6 charge_pump1_0/in5
+ charge_pump1_0/in4 charge_pump1_0/in2 charge_pump1_0/vin m2_6586_52# charge_pump1_0/in8
+ charge_pump1_0/m1_12464_n576# charge_pump1_0/in7 charge_pump1_0/vdd charge_pump1_0/in1
+ VSUBS
Xsky130_fd_pr__nfet_01v8_HRDN5X_0 charge_pump1_0/vdd VSUBS charge_pump1_0/vdd charge_pump1_0/vdd
+ charge_pump1_0/vdd charge_pump1_0/vdd VSUBS VSUBS VSUBS charge_pump1_0/vdd VSUBS
+ charge_pump1_0/vdd VSUBS VSUBS VSUBS VSUBS charge_pump1_0/vdd charge_pump1_0/vdd
+ VSUBS VSUBS VSUBS charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd
+ charge_pump1_0/vdd VSUBS VSUBS VSUBS VSUBS charge_pump1_0/vdd VSUBS sky130_fd_pr__nfet_01v8_HRDN5X
Xcharge_pump1_0 charge_pump1_0/clk_in charge_pump1_0/input1 charge_pump1_0/input2
+ charge_pump1_0/in1 charge_pump1_0/in5 charge_pump1_0/in6 charge_pump1_0/in8 charge_pump1_0/g1
+ charge_pump1_0/g2 charge_pump1_0/clk charge_pump1_0/clkb charge_pump1_0/m1_12464_n576#
+ VSUBS charge_pump1_0/in4 charge_pump1_0/in3 charge_pump1_0/vin charge_pump1_0/vdd
+ charge_pump1_0/in7 charge_pump1_0/in2 VSUBS charge_pump1
Xsky130_fd_pr__nfet_01v8_TKGCLY_0 charge_pump1_0/vdd VSUBS VSUBS VSUBS charge_pump1_0/vdd
+ charge_pump1_0/vdd VSUBS charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd
+ VSUBS VSUBS charge_pump1_0/vdd VSUBS charge_pump1_0/vdd charge_pump1_0/vdd VSUBS
+ VSUBS VSUBS VSUBS charge_pump1_0/vdd VSUBS VSUBS charge_pump1_0/vdd VSUBS charge_pump1_0/vdd
+ charge_pump1_0/vdd charge_pump1_0/vdd VSUBS VSUBS VSUBS VSUBS charge_pump1_0/vdd
+ charge_pump1_0/vdd VSUBS charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd
+ charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd VSUBS
+ VSUBS VSUBS charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd VSUBS VSUBS
+ charge_pump1_0/vdd VSUBS charge_pump1_0/vdd VSUBS VSUBS charge_pump1_0/vdd charge_pump1_0/vdd
+ VSUBS charge_pump1_0/vdd charge_pump1_0/vdd VSUBS VSUBS charge_pump1_0/vdd VSUBS
+ VSUBS charge_pump1_0/vdd VSUBS VSUBS charge_pump1_0/vdd VSUBS VSUBS charge_pump1_0/vdd
+ charge_pump1_0/vdd charge_pump1_0/vdd VSUBS VSUBS VSUBS charge_pump1_0/vdd VSUBS
+ VSUBS VSUBS VSUBS charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd
+ VSUBS VSUBS charge_pump1_0/vdd VSUBS charge_pump1_0/vdd VSUBS charge_pump1_0/vdd
+ VSUBS charge_pump1_0/vdd VSUBS charge_pump1_0/vdd charge_pump1_0/vdd charge_pump1_0/vdd
+ VSUBS VSUBS VSUBS sky130_fd_pr__nfet_01v8_TKGCLY
Xbuffer_digital_0 charge_pump1_0/clk_in m1_7772_199# VSUBS charge_pump1_0/vdd buffer_digital
Xbuffer_digital_1 m1_7772_199# m2_6586_52# VSUBS charge_pump1_0/vdd buffer_digital
Xnmos_decap_10_0 charge_pump1_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_1 charge_pump1_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_2 charge_pump1_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_3 charge_pump1_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_4 charge_pump1_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_6 charge_pump1_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_5 charge_pump1_0/vdd VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_0 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_1 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_2 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_3 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_4 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_5 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_6 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_7 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_9 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_8 VSUBS charge_pump1_0/vdd VSUBS pmos_decap_10
C0 charge_pump1_0/vdd charge_pump1_0/clk_in 5.29f
C1 charge_pump1_0/vdd VSUBS 19.3f
C2 VSUBS m2_6586_52# 3.79f
C3 VSUBS charge_pump1_0/clk_in 9.58f
C4 m2_6586_52# 0 2.92f
C5 charge_pump1_0/input1 0 22.5f
C6 charge_pump1_0/input2 0 22.2f
C7 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C8 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C9 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C10 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C11 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C12 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C13 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C14 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C15 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C16 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C17 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C18 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C19 charge_pump1_0/m1_4341_n519# 0 3.77f
C20 charge_pump1_0/m1_12659_300# 0 2.54f
C21 charge_pump1_0/m1_12464_n576# 0 4.25f
C22 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C23 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C24 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C25 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C26 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C27 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C28 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C29 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C30 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C31 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C32 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C33 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C34 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C35 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C36 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C37 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C38 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C39 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C40 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C41 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C42 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C43 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C44 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C45 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C46 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C47 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C48 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C49 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C50 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C51 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C52 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C53 charge_pump1_0/clkb 0 85.9f
C54 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C55 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C56 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C57 charge_pump1_0/clk 0 85.1f
C58 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C59 charge_pump1_0/vdd 0 0.535p
C60 VSUBS 0 82.2f
C61 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C62 charge_pump1_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C63 charge_pump1_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C64 charge_pump1_0/clock_0/a_344_102# 0 2.81f
C65 charge_pump1_0/clock_0/a_2402_572# 0 2.17f
C66 charge_pump1_0/clock_0/a_344_n986# 0 2.38f
C67 charge_pump1_0/clk_in 0 3.55f
C68 charge_pump1_0/clock_0/a_3246_118# 0 6.83f
C69 charge_pump1_0/g2 0 2.34f
C70 charge_pump1_0/vin 0 10.4f
.ends

.subckt charge_pump1_reverse input1 input2 in1 in5 in6 in8 vdd gnd m1_12464_n576#
+ clock_1/clk_in a_3340_18086# in4 in3 nmos_dnw3_0/vs in7 in2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 nmos_dnw3_0/vs input1 input2 nmos_dnw3_0/clk nmos_dnw3_0/clkb nmos_dnw3_0/vs
+ gnd nmos_dnw3
Xclock_1 clock_1/clk_in vdd gnd clock_1/clk clock_1/clkb clock
Xcapacitor_8_0 vdd input1 vdd clock_1/clkb vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 vdd clock_1/clk vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 in1 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_1 input2 in1 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_2 input1 in2 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 in3 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_4 input2 in2 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_5 input2 in3 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_6 input1 in4 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_7 input1 in5 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_8 input1 in6 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_9 input1 in7 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 in7 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_11 input2 in6 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 in4 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_12 input2 in5 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clock_1/clk input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clock_1/clkb input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 clock_1/clk gnd 2.15f
C1 nmos_dnw3_0/vs clock_1/clkb 2.22f
C2 m1_12464_n576# clock_1/clk 2.14f
C3 vdd clock_1/clk 28.7f
C4 input2 gnd 8.36f
C5 vdd gnd 0.171p
C6 input2 vdd 26.5f
C7 nmos_dnw3_0/vs vdd 9.24f
C8 input1 gnd 8.6f
C9 input2 input1 3.06f
C10 clock_1/clkb gnd 3.21f
C11 input1 vdd 26.5f
C12 m1_12464_n576# clock_1/clkb 2.3f
C13 vdd clock_1/clkb 32.3f
C14 input1 0 22.6f
C15 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C16 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C17 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C18 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C19 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C20 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C21 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C22 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C23 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C24 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C25 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C26 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C27 m1_4341_n519# 0 3.33f
C28 input2 0 22.2f
C29 m1_12659_300# 0 2.68f
C30 m1_12464_n576# 0 4.64f
C31 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C32 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C33 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C34 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C35 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C36 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C37 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C38 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C39 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C40 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C41 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C42 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C43 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C44 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C45 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C46 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C47 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C48 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C49 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C50 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C51 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C52 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C53 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C54 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C55 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C56 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C57 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C58 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C59 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C60 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C61 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C62 clock_1/clk 0 90.7f
C63 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C64 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C65 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C66 clock_1/clkb 0 97.4f
C67 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C68 vdd 0 0.463p
C69 gnd 0 44.4f
C70 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C71 clock_1/a_2432_n962# 0 8.68f **FLOATING
C72 clock_1/a_2020_n482# 0 2.57f **FLOATING
C73 clock_1/a_344_102# 0 2.81f
C74 clock_1/a_2402_572# 0 2.17f
C75 clock_1/a_344_n986# 0 2.38f
C76 clock_1/a_3246_118# 0 6.83f
C77 nmos_dnw3_0/vs 0 10.4f
.ends

.subckt cp1_buffer1_reverse charge_pump1_reverse_0/m1_12464_n576# charge_pump1_reverse_0/in5
+ charge_pump1_reverse_0/clock_1/clk_in charge_pump1_reverse_0/vdd charge_pump1_reverse_0/in8
+ charge_pump1_reverse_0/nmos_dnw3_0/vs charge_pump1_reverse_0/in6 charge_pump1_reverse_0/in1
+ charge_pump1_reverse_0/in4 charge_pump1_reverse_0/in3 m2_6586_52# VSUBS charge_pump1_reverse_0/in7
+ charge_pump1_reverse_0/in2
Xpmos_decap_10_10 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_11 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_12 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_13 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_14 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xcharge_pump1_reverse_0 charge_pump1_reverse_0/input1 charge_pump1_reverse_0/input2
+ charge_pump1_reverse_0/in1 charge_pump1_reverse_0/in5 charge_pump1_reverse_0/in6
+ charge_pump1_reverse_0/in8 charge_pump1_reverse_0/vdd VSUBS charge_pump1_reverse_0/m1_12464_n576#
+ charge_pump1_reverse_0/clock_1/clk_in VSUBS charge_pump1_reverse_0/in4 charge_pump1_reverse_0/in3
+ charge_pump1_reverse_0/nmos_dnw3_0/vs charge_pump1_reverse_0/in7 charge_pump1_reverse_0/in2
+ charge_pump1_reverse
Xbuffer_digital_0 charge_pump1_reverse_0/clock_1/clk_in m1_7766_199# VSUBS charge_pump1_reverse_0/vdd
+ buffer_digital
Xbuffer_digital_1 m1_7766_199# m2_6586_52# VSUBS charge_pump1_reverse_0/vdd buffer_digital
Xnmos_decap_10_0 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_1 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_2 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_3 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_4 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_10 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_11 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_6 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_5 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_12 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_7 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_8 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_0 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xnmos_decap_10_9 charge_pump1_reverse_0/vdd VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_1 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_2 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_3 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_4 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_5 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_6 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_7 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_9 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
Xpmos_decap_10_8 VSUBS charge_pump1_reverse_0/vdd VSUBS pmos_decap_10
C0 VSUBS charge_pump1_reverse_0/vdd 20.3f
C1 charge_pump1_reverse_0/vdd charge_pump1_reverse_0/clock_1/clk_in 5.98f
C2 VSUBS charge_pump1_reverse_0/clock_1/clk_in 12.5f
C3 VSUBS m2_6586_52# 4.22f
C4 charge_pump1_reverse_0/clock_1/clkb charge_pump1_reverse_0/vdd 2.74f
C5 m2_6586_52# 0 2.44f
C6 charge_pump1_reverse_0/input1 0 22.6f
C7 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C8 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C9 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C10 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C11 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C12 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C13 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C14 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C15 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C16 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C17 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C18 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C19 charge_pump1_reverse_0/m1_4341_n519# 0 3.33f
C20 charge_pump1_reverse_0/input2 0 22.2f
C21 charge_pump1_reverse_0/m1_12659_300# 0 2.68f
C22 charge_pump1_reverse_0/m1_12464_n576# 0 4.64f
C23 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C24 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C25 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C26 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C27 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C28 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C29 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C30 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C31 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C32 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C33 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C34 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C35 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C36 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C37 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C38 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C39 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C40 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C41 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C42 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C43 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C44 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C45 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C46 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C47 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C48 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C49 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C50 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C51 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C52 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C53 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C54 charge_pump1_reverse_0/clock_1/clk 0 90.7f
C55 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C56 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C57 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C58 charge_pump1_reverse_0/clock_1/clkb 0 97.4f
C59 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C60 charge_pump1_reverse_0/vdd 0 0.528p
C61 VSUBS 0 87.7f
C62 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C63 charge_pump1_reverse_0/clock_1/a_2432_n962# 0 8.68f **FLOATING
C64 charge_pump1_reverse_0/clock_1/a_2020_n482# 0 2.57f **FLOATING
C65 charge_pump1_reverse_0/clock_1/a_344_102# 0 2.81f
C66 charge_pump1_reverse_0/clock_1/a_2402_572# 0 2.17f
C67 charge_pump1_reverse_0/clock_1/a_344_n986# 0 2.38f
C68 charge_pump1_reverse_0/clock_1/clk_in 0 4f
C69 charge_pump1_reverse_0/clock_1/a_3246_118# 0 6.83f
C70 charge_pump1_reverse_0/nmos_dnw3_0/vs 0 10.4f
.ends

.subckt cp1_buffer_5stage
Xcp1_buffer1_0 cp1_buffer1_0/charge_pump1_0/clk_in cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in4
+ cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_0/charge_pump1_0/vin cp1_buffer1_0/m2_6586_52#
+ cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_2/charge_pump1_0/in7 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in1
+ VSUBS cp1_buffer1
Xcp1_buffer1_1 cp1_buffer1_1/charge_pump1_0/clk_in cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in4
+ cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_1/charge_pump1_0/vin cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in
+ cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_2/charge_pump1_0/in7 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in1
+ VSUBS cp1_buffer1
Xcp1_buffer1_2 cp1_buffer1_2/charge_pump1_0/clk_in cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in4
+ cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/vin cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in
+ cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/m1_12464_n576# cp1_buffer1_2/charge_pump1_0/in7
+ cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in1 VSUBS cp1_buffer1
Xcp1_buffer1_reverse_0 cp1_buffer1_1/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/in4
+ cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_2/charge_pump1_0/vdd
+ cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/in5
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_0/charge_pump1_0/clk_in VSUBS cp1_buffer1_2/charge_pump1_0/in2
+ cp1_buffer1_2/charge_pump1_0/in7 cp1_buffer1_reverse
Xcp1_buffer1_reverse_1 cp1_buffer1_2/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/in4
+ cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_2/charge_pump1_0/vdd
+ cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/in5
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_1/charge_pump1_0/clk_in VSUBS cp1_buffer1_2/charge_pump1_0/in2
+ cp1_buffer1_2/charge_pump1_0/in7 cp1_buffer1_reverse
C0 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in4 3.95f
C1 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in3 3.9f
C2 VSUBS cp1_buffer1_2/charge_pump1_0/in7 3.87f
C3 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in8 3.7f
C4 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/vdd 3.91f
C5 VSUBS cp1_buffer1_0/charge_pump1_0/clk_in 3.12f
C6 VSUBS cp1_buffer1_2/charge_pump1_0/in6 4.33f
C7 cp1_buffer1_2/charge_pump1_0/vdd VSUBS 79.4f
C8 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in2 3.97f
C9 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in1 4f
C10 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in 4.13f
C11 VSUBS cp1_buffer1_2/charge_pump1_0/in4 4.19f
C12 VSUBS cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in 2.12f
C13 VSUBS cp1_buffer1_2/charge_pump1_0/in3 4.13f
C14 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/clk_in 2.55f
C15 VSUBS cp1_buffer1_2/charge_pump1_0/in8 3.81f
C16 cp1_buffer1_2/charge_pump1_0/in5 VSUBS 4.13f
C17 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in7 3.64f
C18 VSUBS cp1_buffer1_2/charge_pump1_0/in2 4.24f
C19 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/clk_in 2.01f
C20 VSUBS cp1_buffer1_2/charge_pump1_0/in1 4.13f
C21 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in6 4.05f
C22 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in VSUBS 2.14f
C23 VSUBS cp1_buffer1_1/charge_pump1_0/clk_in 3.35f
C24 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 0 22.6f
C25 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C26 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C27 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C28 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C29 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C30 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C31 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C32 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C33 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C34 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C35 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C36 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C37 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_4341_n519# 0 3.33f
C38 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 0 22.2f
C39 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_12659_300# 0 2.68f
C40 cp1_buffer1_2/charge_pump1_0/vin 0 13.3f
C41 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C42 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C43 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C44 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C45 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C46 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C47 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C48 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C49 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C50 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C51 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C52 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C53 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C54 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C55 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C56 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C57 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C58 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C59 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C60 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C61 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C62 cp1_buffer1_2/charge_pump1_0/in6 0 7.43f
C63 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C64 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C65 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C66 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C67 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C68 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C69 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C70 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C71 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C72 cp1_buffer1_2/charge_pump1_0/in8 0 7.77f
C73 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C74 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk 0 90.7f
C75 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C76 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C77 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C78 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb 0 97.4f
C79 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C80 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C81 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2432_n962# 0 8.68f **FLOATING
C82 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2020_n482# 0 2.57f **FLOATING
C83 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_102# 0 2.81f
C84 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2402_572# 0 2.17f
C85 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_n986# 0 2.38f
C86 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in 0 7.19f
C87 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_3246_118# 0 6.83f
C88 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 0 22.6f
C89 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C90 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C91 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C92 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C93 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C94 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C95 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C96 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C97 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C98 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C99 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C100 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C101 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_4341_n519# 0 3.33f
C102 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 0 22.2f
C103 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_12659_300# 0 2.68f
C104 cp1_buffer1_1/charge_pump1_0/vin 0 13.2f
C105 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C106 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C107 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C108 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C109 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C110 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C111 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C112 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C113 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C114 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C115 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C116 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C117 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C118 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C119 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C120 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C121 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C122 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C123 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C124 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C125 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C126 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C127 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C128 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C129 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C130 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C131 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C132 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C133 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C134 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C135 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C136 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 0 90.7f
C137 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C138 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C139 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C140 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb 0 97.4f
C141 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C142 cp1_buffer1_2/charge_pump1_0/vdd 0 2.67p
C143 VSUBS 0 0.421p
C144 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C145 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2432_n962# 0 8.68f **FLOATING
C146 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2020_n482# 0 2.57f **FLOATING
C147 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_102# 0 2.81f
C148 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2402_572# 0 2.17f
C149 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_n986# 0 2.38f
C150 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in 0 5.18f
C151 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_3246_118# 0 6.83f
C152 cp1_buffer1_2/charge_pump1_0/input1 0 22.5f
C153 cp1_buffer1_2/charge_pump1_0/input2 0 22.2f
C154 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C155 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C156 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C157 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C158 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C159 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C160 cp1_buffer1_2/charge_pump1_0/in4 0 7.51f
C161 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C162 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C163 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C164 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C165 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C166 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C167 cp1_buffer1_2/charge_pump1_0/m1_4341_n519# 0 3.77f
C168 cp1_buffer1_2/charge_pump1_0/m1_12659_300# 0 2.54f
C169 cp1_buffer1_2/charge_pump1_0/m1_12464_n576# 0 4.25f
C170 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C171 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C172 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C173 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C174 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C175 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C176 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C177 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C178 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C179 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C180 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C181 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C182 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C183 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C184 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C185 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C186 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C187 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C188 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C189 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C190 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C191 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C192 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C193 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C194 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C195 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C196 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C197 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C198 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C199 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C200 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C201 cp1_buffer1_2/charge_pump1_0/clkb 0 85.9f
C202 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C203 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C204 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C205 cp1_buffer1_2/charge_pump1_0/clk 0 85.1f
C206 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C207 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C208 cp1_buffer1_2/charge_pump1_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C209 cp1_buffer1_2/charge_pump1_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C210 cp1_buffer1_2/charge_pump1_0/clock_0/a_344_102# 0 2.81f
C211 cp1_buffer1_2/charge_pump1_0/clock_0/a_2402_572# 0 2.17f
C212 cp1_buffer1_2/charge_pump1_0/clock_0/a_344_n986# 0 2.38f
C213 cp1_buffer1_2/charge_pump1_0/clk_in 0 3.55f
C214 cp1_buffer1_2/charge_pump1_0/clock_0/a_3246_118# 0 6.83f
C215 cp1_buffer1_2/charge_pump1_0/g2 0 2.34f
C216 cp1_buffer1_1/charge_pump1_0/input1 0 22.5f
C217 cp1_buffer1_1/charge_pump1_0/input2 0 22.2f
C218 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C219 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C220 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C221 cp1_buffer1_2/charge_pump1_0/in5 0 7.49f
C222 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C223 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C224 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C225 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C226 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C227 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C228 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C229 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C230 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C231 cp1_buffer1_1/charge_pump1_0/m1_4341_n519# 0 3.77f
C232 cp1_buffer1_1/charge_pump1_0/m1_12659_300# 0 2.54f
C233 cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs 0 14.5f
C234 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C235 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C236 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C237 cp1_buffer1_2/charge_pump1_0/in7 0 7.35f
C238 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C239 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C240 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C241 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C242 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C243 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C244 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C245 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C246 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C247 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C248 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C249 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C250 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C251 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C252 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C253 cp1_buffer1_2/charge_pump1_0/in2 0 7.41f
C254 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C255 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C256 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C257 cp1_buffer1_2/charge_pump1_0/in3 0 7.39f
C258 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C259 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C260 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C261 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C262 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C263 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C264 cp1_buffer1_2/charge_pump1_0/in1 0 7.1f
C265 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C266 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C267 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C268 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C269 cp1_buffer1_1/charge_pump1_0/clkb 0 85.9f
C270 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C271 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C272 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C273 cp1_buffer1_1/charge_pump1_0/clk 0 85.1f
C274 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C275 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C276 cp1_buffer1_1/charge_pump1_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C277 cp1_buffer1_1/charge_pump1_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C278 cp1_buffer1_1/charge_pump1_0/clock_0/a_344_102# 0 2.81f
C279 cp1_buffer1_1/charge_pump1_0/clock_0/a_2402_572# 0 2.17f
C280 cp1_buffer1_1/charge_pump1_0/clock_0/a_344_n986# 0 2.38f
C281 cp1_buffer1_1/charge_pump1_0/clock_0/a_3246_118# 0 6.83f
C282 cp1_buffer1_1/charge_pump1_0/g2 0 2.34f
C283 cp1_buffer1_0/m2_6586_52# 0 2.92f
C284 cp1_buffer1_0/charge_pump1_0/input1 0 22.5f
C285 cp1_buffer1_0/charge_pump1_0/input2 0 22.2f
C286 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C287 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C288 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C289 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C290 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C291 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C292 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C293 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C294 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C295 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C296 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C297 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C298 cp1_buffer1_0/charge_pump1_0/m1_4341_n519# 0 3.77f
C299 cp1_buffer1_0/charge_pump1_0/m1_12659_300# 0 2.54f
C300 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs 0 14.6f
C301 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C302 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C303 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C304 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C305 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C306 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C307 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C308 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C309 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C310 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C311 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C312 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C313 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C314 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C315 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C316 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C317 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C318 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C319 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C320 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C321 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C322 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C323 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C324 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C325 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C326 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C327 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C328 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C329 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C330 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C331 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C332 cp1_buffer1_0/charge_pump1_0/clkb 0 85.9f
C333 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C334 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C335 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C336 cp1_buffer1_0/charge_pump1_0/clk 0 85.1f
C337 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C338 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C339 cp1_buffer1_0/charge_pump1_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C340 cp1_buffer1_0/charge_pump1_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C341 cp1_buffer1_0/charge_pump1_0/clock_0/a_344_102# 0 2.81f
C342 cp1_buffer1_0/charge_pump1_0/clock_0/a_2402_572# 0 2.17f
C343 cp1_buffer1_0/charge_pump1_0/clock_0/a_344_n986# 0 2.38f
C344 cp1_buffer1_0/charge_pump1_0/clk_in 0 3.27f
C345 cp1_buffer1_0/charge_pump1_0/clock_0/a_3246_118# 0 6.83f
C346 cp1_buffer1_0/charge_pump1_0/g2 0 2.34f
C347 cp1_buffer1_0/charge_pump1_0/vin 0 10.4f
.ends

