magic
tech sky130A
magscale 1 2
timestamp 1698861456
<< locali >>
rect 2418 3468 4121 3477
rect 2418 3430 3518 3431
rect 2418 3409 2604 3430
rect 2672 3300 2742 3428
rect 2876 3409 3518 3430
rect 3598 3409 4121 3431
rect 3836 3304 3900 3409
rect 4840 3362 5016 3396
rect 2806 3218 2890 3220
rect 3658 3218 3964 3224
rect 2806 3217 3034 3218
rect 2634 3176 3034 3217
rect 3544 3176 3964 3218
rect 3658 3169 3964 3176
rect 3658 3168 3730 3169
rect 3894 3166 3964 3169
rect 2678 2752 2746 2888
rect 3834 2748 3902 2888
rect 2506 2636 2810 2704
rect 3662 2620 3970 2704
rect 4843 2665 4864 2747
rect 5047 2596 5129 2606
rect 4369 2494 4451 2496
rect 5047 2494 5129 2496
rect 3234 2486 5376 2494
rect 3146 2484 5376 2486
rect 2420 2474 5376 2484
rect 2420 2428 5018 2437
rect 5363 2437 5376 2474
rect 5134 2428 5376 2437
rect 2420 2426 4158 2428
<< viali >>
rect 2415 3434 4123 3468
rect 2415 3431 3518 3434
rect 3598 3431 4123 3434
rect 2414 2438 5363 2474
rect 2414 2437 5018 2438
rect 5134 2437 5363 2438
<< metal1 >>
rect 4954 3526 4964 3584
rect 5156 3526 5166 3584
rect 4984 3522 5157 3526
rect 2418 3474 4121 3477
rect 2403 3468 4135 3474
rect 2403 3431 2415 3468
rect 3518 3431 3598 3434
rect 4123 3431 4135 3468
rect 2403 3425 4135 3431
rect 2418 3410 4121 3425
rect 2418 3409 3518 3410
rect 3598 3409 4121 3410
rect 2598 3408 2916 3409
rect 2971 3408 3010 3409
rect 3737 3406 3775 3409
rect 4984 3396 5156 3421
rect 4881 3362 5156 3396
rect 3146 3158 3250 3216
rect 2976 3110 3180 3120
rect 2976 3058 2992 3110
rect 3168 3058 3180 3110
rect 2976 3044 3180 3058
rect 3212 2718 3250 3158
rect 3307 3177 3410 3216
rect 3307 2720 3346 3177
rect 3396 3108 3600 3114
rect 3396 3046 3406 3108
rect 3578 3046 3600 3108
rect 4881 3073 4915 3362
rect 4984 3342 5156 3362
rect 4948 3200 4958 3258
rect 5150 3200 5160 3258
rect 4984 3073 5158 3104
rect 3396 3038 3600 3046
rect 4879 3039 5158 3073
rect 4879 2761 4913 3039
rect 4984 3025 5158 3039
rect 4942 2880 4952 2938
rect 5144 2880 5154 2938
rect 4984 2761 5158 2785
rect 4879 2727 5158 2761
rect 1624 2482 1634 2686
rect 2102 2482 2112 2686
rect 2972 2616 2982 2707
rect 3039 2616 3049 2707
rect 3182 2703 3250 2718
rect 3306 2708 3424 2720
rect 3148 2702 3250 2703
rect 3136 2616 3146 2702
rect 3204 2628 3250 2702
rect 3204 2616 3222 2628
rect 3302 2616 3312 2708
rect 3422 2616 3432 2708
rect 3532 2642 3542 2714
rect 3596 2642 3606 2714
rect 4984 2706 5158 2727
rect 3148 2614 3222 2616
rect 3306 2614 3319 2616
rect 3392 2614 3424 2616
rect 3306 2612 3424 2614
rect 4948 2564 4958 2622
rect 5150 2564 5160 2622
rect 5204 2614 5245 3501
rect 4984 2562 5036 2564
rect 3234 2494 3510 2495
rect 3958 2494 4121 2495
rect 3234 2486 5376 2494
rect 3146 2484 5376 2486
rect 2396 2474 5376 2484
rect 2396 2437 2414 2474
rect 5018 2437 5134 2438
rect 5363 2437 5376 2474
rect 2396 2428 5376 2437
rect 2396 2427 4158 2428
rect 2396 2424 2430 2427
rect 4090 2426 4158 2427
rect 5500 2418 5506 2532
rect 5496 436 5506 2418
rect 5626 436 5636 2532
<< via1 >>
rect 4964 3526 5156 3584
rect 2992 3058 3168 3110
rect 3406 3046 3578 3108
rect 4958 3200 5150 3258
rect 4952 2880 5144 2938
rect 1634 2482 2102 2686
rect 2982 2616 3039 2707
rect 3146 2616 3204 2702
rect 3312 2616 3422 2708
rect 3542 2642 3596 2714
rect 3319 2614 3392 2616
rect 4958 2564 5150 2622
rect 5506 436 5626 2532
<< metal2 >>
rect 4948 3584 5160 3598
rect 4948 3526 4964 3584
rect 5156 3526 5160 3584
rect 4948 3258 5160 3526
rect 4948 3200 4958 3258
rect 5150 3200 5160 3258
rect 2976 3114 3180 3120
rect 3406 3114 3578 3118
rect 2976 3110 3600 3114
rect 2976 3058 2992 3110
rect 3168 3108 3600 3110
rect 3168 3076 3406 3108
rect 3168 3058 3180 3076
rect 2976 3044 3180 3058
rect 3396 3046 3406 3076
rect 3578 3046 3600 3108
rect 3396 3038 3600 3046
rect 3406 3036 3578 3038
rect 4948 2967 5160 3200
rect 3000 2938 5160 2967
rect 3000 2928 4952 2938
rect 3000 2717 3039 2928
rect 3544 2724 3583 2928
rect 4948 2880 4952 2928
rect 5144 2880 5160 2938
rect 2982 2707 3039 2717
rect 1634 2686 2102 2696
rect 2982 2610 3039 2616
rect 3146 2702 3204 2712
rect 3146 2610 3204 2616
rect 3306 2708 3424 2720
rect 3306 2616 3312 2708
rect 3422 2616 3424 2708
rect 3542 2714 3596 2724
rect 3596 2646 3598 2696
rect 3542 2632 3596 2642
rect 3544 2630 3583 2632
rect 3306 2614 3319 2616
rect 3392 2614 3424 2616
rect 3306 2612 3424 2614
rect 4948 2622 5160 2880
rect 2102 2578 2342 2580
rect 3156 2578 3204 2610
rect 2102 2576 3204 2578
rect 3307 2606 3422 2612
rect 2102 2496 3206 2576
rect 2102 2494 2324 2496
rect 2352 2494 2412 2496
rect 2102 2484 2134 2494
rect 1634 2472 2102 2482
rect 3307 2416 3348 2606
rect 4948 2564 4958 2622
rect 5150 2564 5160 2622
rect 4948 2556 5160 2564
rect 4958 2554 5150 2556
rect 5506 2532 5626 2542
rect 5500 2489 5506 2530
rect 3307 2375 5506 2416
rect 3307 2372 3348 2375
rect 5506 426 5626 436
<< via2 >>
rect 1648 2496 2064 2666
rect 5506 436 5626 2532
<< metal3 >>
rect 1608 2472 1618 2702
rect 2120 2472 2130 2702
rect 5500 2532 5636 2537
rect 5500 2423 5506 2532
rect 5496 436 5506 2423
rect 5626 436 5636 2532
rect 5496 431 5636 436
<< via3 >>
rect 1618 2666 2120 2702
rect 1618 2496 1648 2666
rect 1648 2496 2064 2666
rect 2064 2496 2120 2666
rect 1618 2472 2120 2496
<< metal4 >>
rect 1617 2702 2121 2703
rect 1617 2472 1618 2702
rect 2120 2472 2121 2702
rect 1617 2471 2121 2472
rect 1682 1960 1934 2471
use sky130_fd_pr__nfet_01v8_EJYG4R  sky130_fd_pr__nfet_01v8_EJYG4R_0
timestamp 1697915631
transform 0 -1 5088 1 0 3064
box -641 -279 641 279
use sky130_fd_pr__nfet_01v8_SMGLWN  sky130_fd_pr__nfet_01v8_SMGLWN_0
timestamp 1698155087
transform 1 0 2712 0 1 2667
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  sky130_fd_pr__nfet_01v8_SMGLWN_1
timestamp 1698155087
transform 1 0 3870 0 1 2667
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_lvt_TM5SY6  sky130_fd_pr__pfet_01v8_lvt_TM5SY6_0
timestamp 1698622305
transform 1 0 3868 0 1 3208
box -246 -269 246 269
use sky130_fd_pr__cap_mim_m3_1_TNHPNJ  XC3
timestamp 1697379271
transform 1 0 3433 0 1 1299
box -2186 -1040 2186 1040
use sky130_fd_pr__nfet_01v8_SMGLWN  XM1
timestamp 1698155087
transform 1 0 3098 0 1 2667
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM2
timestamp 1698155087
transform 1 0 3484 0 1 2667
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_lvt_TM5SY6  XM3
timestamp 1698622305
transform 1 0 3482 0 1 3208
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_lvt_TM5SY6  XM6
timestamp 1698622305
transform 1 0 2710 0 1 3208
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_lvt_TM5SY6  XM18
timestamp 1698622305
transform 1 0 3096 0 1 3208
box -246 -269 246 269
<< labels >>
rlabel metal2 4602 2416 4602 2416 1 vo1
rlabel viali 4134 2455 4134 2455 3 gnd
rlabel metal1 4056 3477 4056 3477 1 Vdd
<< end >>
