magic
tech sky130A
magscale 1 2
timestamp 1698329102
<< nwell >>
rect 4998 -7520 5006 -6164
rect 4998 -7526 5272 -7520
<< psubdiff >>
rect -2060 -6652 1008 -6518
rect -2060 -7070 -1906 -6652
rect 796 -7070 1008 -6652
rect -2060 -7208 1008 -7070
rect 11210 -6708 14266 -6598
rect 11210 -7178 11356 -6708
rect 14084 -7178 14266 -6708
rect 11210 -7274 14266 -7178
rect 5700 -25120 5830 -25098
rect 5700 -25358 5732 -25120
rect 5796 -25358 5830 -25120
rect 5700 -25384 5830 -25358
<< nsubdiff >>
rect 5038 -7124 5136 -7098
rect 5038 -7418 5064 -7124
rect 5108 -7418 5136 -7124
rect 5038 -7446 5136 -7418
rect 5702 -24868 5828 -24854
rect 5702 -24924 5728 -24868
rect 5790 -24924 5828 -24868
rect 5702 -24944 5828 -24924
<< psubdiffcont >>
rect -1906 -7070 796 -6652
rect 11356 -7178 14084 -6708
rect 5732 -25358 5796 -25120
<< nsubdiffcont >>
rect 5064 -7418 5108 -7124
rect 5728 -24924 5790 -24868
<< poly >>
rect 5324 -6246 5540 -6236
rect 5324 -6288 5358 -6246
rect 5516 -6288 5540 -6246
rect 5324 -6306 5540 -6288
rect 5510 -6460 5540 -6306
rect 6098 -6288 6328 -6272
rect 6098 -6328 6150 -6288
rect 6304 -6328 6328 -6288
rect 6098 -6342 6328 -6328
rect 6098 -6462 6128 -6342
<< polycont >>
rect 5358 -6288 5516 -6246
rect 6150 -6328 6304 -6288
<< locali >>
rect 5322 -6246 5540 -6240
rect 5322 -6288 5358 -6246
rect 5516 -6288 5540 -6246
rect 5322 -6296 5540 -6288
rect 6130 -6288 6328 -6272
rect 6130 -6328 6150 -6288
rect 6304 -6328 6328 -6288
rect 6130 -6342 6328 -6328
rect -2060 -6652 1008 -6518
rect -2060 -7070 -1906 -6652
rect 796 -7070 1008 -6652
rect -2060 -7208 1008 -7070
rect 11210 -6708 14266 -6598
rect 5038 -7124 5136 -7098
rect 5038 -7418 5064 -7124
rect 5108 -7418 5136 -7124
rect 11210 -7178 11356 -6708
rect 14084 -7178 14266 -6708
rect 11210 -7274 14266 -7178
rect 5038 -7446 5136 -7418
rect 5702 -24868 5828 -24854
rect 5702 -24924 5728 -24868
rect 5790 -24924 5828 -24868
rect 5702 -24944 5828 -24924
rect 5700 -25120 5830 -25098
rect 5700 -25358 5732 -25120
rect 5796 -25358 5830 -25120
rect 5700 -25384 5830 -25358
<< viali >>
rect 5358 -6288 5516 -6246
rect 6150 -6328 6304 -6288
rect -1906 -7070 796 -6652
rect 5064 -7418 5108 -7124
rect 11356 -7178 14084 -6708
rect 5728 -24924 5790 -24868
rect 5732 -25358 5796 -25120
<< metal1 >>
rect 5322 -6294 5358 -6240
rect 5516 -6294 5540 -6240
rect 5322 -6296 5540 -6294
rect 6130 -6278 6328 -6272
rect 6130 -6334 6146 -6278
rect 6314 -6334 6328 -6278
rect 6130 -6342 6328 -6334
rect -2060 -6652 1008 -6518
rect 5308 -6556 5502 -6488
rect 6134 -6562 6338 -6488
rect -2060 -7070 -1906 -6652
rect 796 -7070 1008 -6652
rect -2060 -7208 1008 -7070
rect 5046 -7124 5136 -7098
rect 5046 -7371 5064 -7124
rect -4887 -7418 5064 -7371
rect 5108 -7418 5136 -7124
rect 5308 -7208 5424 -6630
rect 6224 -7212 6338 -6634
rect 11210 -6708 14266 -6598
rect 11210 -7178 11356 -6708
rect 14084 -7178 14266 -6708
rect 11210 -7274 14266 -7178
rect -4887 -7434 5136 -7418
rect -4887 -7473 5133 -7434
rect -4887 -24732 -4785 -7473
rect 5312 -7506 5390 -7316
rect 3184 -11121 3413 -11087
rect 3260 -17375 3467 -17341
rect 3258 -23423 3413 -23389
rect 15638 -24730 15834 -24674
rect -4887 -24800 5830 -24732
rect -4887 -24802 -4785 -24800
rect 5700 -24868 5830 -24800
rect 5700 -24924 5728 -24868
rect 5790 -24924 5830 -24868
rect 5564 -25090 5636 -25080
rect -4274 -25622 -4054 -25588
rect -4274 -26806 -4240 -25622
rect -4084 -26806 -4054 -25622
rect 5564 -25668 5576 -25090
rect 5630 -25668 5636 -25090
rect 5700 -25120 5830 -24924
rect 5700 -25358 5732 -25120
rect 5796 -25358 5830 -25120
rect 5700 -25384 5830 -25358
rect 5918 -25088 6004 -25056
rect 5564 -25676 5636 -25668
rect 5918 -25666 5932 -25088
rect 5990 -25666 6004 -25088
rect 5918 -25676 6004 -25666
rect 5750 -25984 5786 -25852
rect -4274 -26819 -4054 -26806
rect 15638 -26798 15672 -24730
rect 15798 -26798 15834 -24730
rect -4274 -26853 5758 -26819
rect 15638 -26820 15834 -26798
rect -4274 -26860 -4054 -26853
rect 5724 -26977 5758 -26853
rect 5864 -26854 15834 -26820
rect 5864 -26856 15758 -26854
rect 5864 -26986 5900 -26856
<< via1 >>
rect 5358 -6246 5516 -6240
rect 5358 -6288 5516 -6246
rect 5358 -6294 5516 -6288
rect 6146 -6288 6314 -6278
rect 6146 -6328 6150 -6288
rect 6150 -6328 6304 -6288
rect 6304 -6328 6314 -6288
rect 6146 -6334 6314 -6328
rect -1906 -7070 796 -6652
rect 11356 -7178 14084 -6708
rect -4240 -26806 -4084 -25622
rect 5576 -25668 5630 -25090
rect 5932 -25666 5990 -25088
rect 15672 -26798 15798 -24730
<< metal2 >>
rect 4672 -6220 4988 -6218
rect 4594 -6236 4988 -6220
rect 4594 -6310 4612 -6236
rect 4964 -6240 4988 -6236
rect 4964 -6294 5358 -6240
rect 5516 -6242 5540 -6240
rect 5516 -6294 6096 -6242
rect 4964 -6296 6096 -6294
rect 4964 -6310 4988 -6296
rect 5296 -6298 6096 -6296
rect 6130 -6276 6328 -6272
rect 6130 -6278 6150 -6276
rect 6304 -6278 6328 -6276
rect 4594 -6324 4988 -6310
rect 4594 -6326 4986 -6324
rect 6130 -6334 6146 -6278
rect 6314 -6334 6328 -6278
rect 6130 -6336 6150 -6334
rect 6304 -6336 6328 -6334
rect 6130 -6342 6328 -6336
rect -2060 -6652 1008 -6518
rect -2060 -7070 -1906 -6652
rect 796 -7070 1008 -6652
rect -2060 -7208 1008 -7070
rect 11210 -6708 14266 -6598
rect 11210 -7178 11356 -6708
rect 14084 -7178 14266 -6708
rect 11210 -7274 14266 -7178
rect 4940 -8782 6692 -8742
rect 4934 -10866 6644 -10826
rect 4962 -12948 6642 -12908
rect 4926 -15034 6600 -14994
rect 4928 -17120 6576 -17080
rect 4934 -19202 6592 -19162
rect 4922 -21290 6656 -21250
rect 4926 -23374 6656 -23334
rect 15638 -24730 15834 -24674
rect 5562 -25090 5644 -25080
rect -4274 -25622 -4054 -25588
rect -4274 -26806 -4240 -25622
rect -4084 -26806 -4054 -25622
rect 5562 -25668 5576 -25090
rect 5632 -25668 5644 -25090
rect 5562 -25676 5644 -25668
rect 5918 -25088 6004 -25056
rect 5918 -25666 5932 -25088
rect 5990 -25666 6004 -25088
rect 5918 -25676 6004 -25666
rect -4274 -26860 -4054 -26806
rect 15638 -26798 15672 -24730
rect 15798 -26798 15834 -24730
rect 15638 -26854 15834 -26798
<< via2 >>
rect 4612 -6310 4964 -6236
rect 6150 -6278 6304 -6276
rect 6150 -6334 6304 -6278
rect 6150 -6336 6304 -6334
rect -1906 -7070 796 -6652
rect 11356 -7178 14084 -6708
rect -4240 -26806 -4084 -25622
rect 5576 -25668 5630 -25090
rect 5630 -25668 5632 -25090
rect 5932 -25666 5990 -25088
rect 15672 -26798 15798 -24730
<< metal3 >>
rect 2360 -6136 4232 -5766
rect -4272 -6345 4232 -6136
rect 7552 -5774 9426 -5766
rect 7552 -6010 9434 -5774
rect 7552 -6202 15831 -6010
rect 4594 -6236 4986 -6218
rect 4594 -6310 4612 -6236
rect 4964 -6310 4986 -6236
rect 4594 -6324 4986 -6310
rect 6132 -6276 6328 -6268
rect 6132 -6336 6150 -6276
rect 6304 -6336 6328 -6276
rect 6132 -6342 6328 -6336
rect 6796 -6276 7268 -6272
rect 6796 -6340 6842 -6276
rect 7246 -6340 7268 -6276
rect 6796 -6342 7268 -6340
rect -4272 -8922 -4063 -6345
rect -2060 -6652 1008 -6518
rect -2060 -7070 -1906 -6652
rect 796 -7070 1008 -6652
rect -2060 -7208 1008 -7070
rect 2360 -7640 4232 -6345
rect 5632 -8846 5744 -7256
rect -4272 -9012 -3980 -8922
rect 4698 -8958 5744 -8846
rect 5912 -8840 6024 -7242
rect 7552 -7636 9434 -6202
rect 11210 -6708 14266 -6598
rect 11210 -7178 11356 -6708
rect 14084 -7178 14266 -6708
rect 11210 -7274 14266 -7178
rect 7552 -7640 9426 -7636
rect 5912 -8952 6852 -8840
rect 15639 -8914 15831 -6202
rect 15584 -8921 15832 -8914
rect 15572 -9003 15832 -8921
rect 15584 -9006 15832 -9003
rect -4272 -11006 -4063 -9012
rect 15639 -11000 15831 -9006
rect -4272 -11098 -3922 -11006
rect 15582 -11090 15831 -11000
rect -4272 -13086 -4063 -11098
rect 15639 -13082 15831 -11090
rect -4272 -13178 -3940 -13086
rect 15586 -13172 15831 -13082
rect -4272 -15170 -4063 -13178
rect 15639 -15168 15831 -13172
rect -4272 -15262 -3916 -15170
rect 15524 -15258 15831 -15168
rect -4272 -17260 -4063 -15262
rect 15639 -17252 15831 -15258
rect -4272 -17352 -3916 -17260
rect 15518 -17342 15831 -17252
rect -4272 -19340 -4063 -17352
rect 15639 -19334 15831 -17342
rect -4272 -19432 -3898 -19340
rect 15512 -19424 15831 -19334
rect -4272 -21428 -4063 -19432
rect 15639 -21424 15831 -19424
rect -4272 -21520 -3898 -21428
rect 15510 -21514 15831 -21424
rect -4272 -23514 -4063 -21520
rect 15639 -23507 15831 -21514
rect -4272 -23597 -3892 -23514
rect 15421 -23589 15831 -23507
rect -4272 -23604 -3896 -23597
rect -4272 -24810 -4063 -23604
rect 1170 -24810 3042 -24562
rect 3398 -24644 4198 -24600
rect 3398 -24770 3440 -24644
rect 4138 -24684 4198 -24644
rect 7200 -24654 7794 -24610
rect 8556 -24636 10428 -24568
rect 5918 -24668 6586 -24656
rect 4138 -24744 5644 -24684
rect 4138 -24770 4198 -24744
rect 3398 -24800 4198 -24770
rect -4272 -25019 3042 -24810
rect -4272 -25588 -4063 -25019
rect -4274 -25622 -4054 -25588
rect -4274 -26806 -4240 -25622
rect -4084 -26806 -4054 -25622
rect 1170 -26430 3042 -25019
rect 5562 -25090 5644 -24744
rect 5562 -25668 5576 -25090
rect 5632 -25668 5644 -25090
rect 5562 -25676 5644 -25668
rect 5918 -24752 7200 -24668
rect 5918 -25056 6002 -24752
rect 7762 -24780 7794 -24654
rect 7200 -24792 7794 -24780
rect 8558 -24758 10428 -24636
rect 15639 -24674 15831 -23589
rect 15638 -24730 15834 -24674
rect 15638 -24758 15672 -24730
rect 8558 -24950 15672 -24758
rect 5918 -25088 6004 -25056
rect 5918 -25666 5932 -25088
rect 5990 -25666 6004 -25088
rect 5918 -25676 6004 -25666
rect 8558 -26440 10428 -24950
rect 8558 -26442 10250 -26440
rect -4274 -26860 -4054 -26806
rect 15638 -26798 15672 -24950
rect 15798 -26798 15834 -24730
rect 15638 -26854 15834 -26798
<< via3 >>
rect 4612 -6310 4964 -6236
rect 6842 -6340 7246 -6276
rect -1906 -7070 796 -6652
rect 11356 -7178 14084 -6708
rect 3440 -24770 4138 -24644
rect 7200 -24780 7762 -24654
<< mimcap >>
rect 2400 -6236 4202 -5798
rect 2400 -6316 3726 -6236
rect 4108 -6316 4202 -6236
rect 2400 -7600 4202 -6316
rect 7600 -6272 9402 -5798
rect 7600 -6338 7670 -6272
rect 7960 -6338 9402 -6272
rect 7600 -7600 9402 -6338
rect 1198 -24634 3002 -24598
rect 1198 -24772 2118 -24634
rect 2874 -24772 3002 -24634
rect 1198 -26400 3002 -24772
rect 8592 -24654 10400 -24598
rect 8592 -24750 8642 -24654
rect 9134 -24750 10400 -24654
rect 8592 -26412 10400 -24750
<< mimcapcontact >>
rect 3726 -6316 4108 -6236
rect 7670 -6338 7960 -6272
rect 2118 -24772 2874 -24634
rect 8642 -24750 9134 -24654
<< metal4 >>
rect 4594 -6220 4986 -6218
rect 3689 -6236 4986 -6220
rect 3689 -6316 3726 -6236
rect 4108 -6310 4612 -6236
rect 4964 -6310 4986 -6236
rect 4108 -6316 4986 -6310
rect 3689 -6324 4986 -6316
rect 6796 -6276 7670 -6272
rect 3689 -6326 4950 -6324
rect 6796 -6340 6842 -6276
rect 7246 -6338 7670 -6276
rect 7960 -6338 7993 -6272
rect 7246 -6340 7993 -6338
rect 6796 -6342 7993 -6340
rect -2060 -6652 1008 -6518
rect -2060 -7070 -1906 -6652
rect 796 -7070 1008 -6652
rect -2060 -7208 1008 -7070
rect 11210 -6708 14266 -6598
rect 11210 -7178 11356 -6708
rect 14084 -7178 14266 -6708
rect 11210 -7274 14266 -7178
rect 15388 -7764 15834 -7762
rect -4934 -8330 -3202 -7774
rect -4934 -9868 -4378 -8330
rect 3462 -8344 8248 -7776
rect 15328 -8331 16459 -7764
rect 15402 -8332 15750 -8331
rect 15892 -9844 16459 -8331
rect -4934 -10424 -3460 -9868
rect 3372 -10416 8158 -9848
rect 15065 -10411 16459 -9844
rect -4934 -11942 -4378 -10424
rect 15892 -11942 16459 -10411
rect -4934 -12496 -3382 -11942
rect -4934 -12498 -4288 -12496
rect -3988 -12498 -3382 -12496
rect -4934 -14014 -4378 -12498
rect 3462 -12528 8248 -11960
rect 15315 -12509 16459 -11942
rect 15892 -14005 16459 -12509
rect -4934 -14568 -3528 -14014
rect -4934 -14570 -4288 -14568
rect -3988 -14570 -3528 -14568
rect -4934 -16126 -4378 -14570
rect 3486 -14596 8424 -14016
rect 15199 -14572 16459 -14005
rect -4934 -16680 -3444 -16126
rect 3334 -16678 8272 -16098
rect 15892 -16104 16459 -14572
rect 15131 -16671 16459 -16104
rect -4934 -16682 -4288 -16680
rect -3988 -16682 -3444 -16680
rect -4934 -18176 -4378 -16682
rect 15892 -18176 16459 -16671
rect -4934 -18182 -3880 -18176
rect -4934 -18732 -3432 -18182
rect -4934 -20282 -4378 -18732
rect 3312 -18768 8250 -18188
rect 15225 -18743 16459 -18176
rect -4934 -20838 -3342 -20282
rect -4934 -22374 -4378 -20838
rect 3428 -20852 8366 -20272
rect 15892 -20274 16459 -18743
rect 15249 -20841 16459 -20274
rect -4934 -22930 -2608 -22374
rect 3440 -22936 8378 -22356
rect 15892 -22364 16459 -20841
rect 15023 -22931 16459 -22364
rect 2048 -24634 4198 -24598
rect 2048 -24772 2118 -24634
rect 2874 -24644 4198 -24634
rect 2874 -24770 3440 -24644
rect 4138 -24770 4198 -24644
rect 2874 -24772 4198 -24770
rect 2048 -24802 4198 -24772
rect 7194 -24654 9202 -24618
rect 7194 -24780 7200 -24654
rect 7762 -24750 8642 -24654
rect 9134 -24750 9202 -24654
rect 7762 -24780 9202 -24750
rect 7194 -24800 9202 -24780
rect 15892 -28844 16459 -22931
rect 7049 -29411 16459 -28844
<< via4 >>
rect -1906 -7070 796 -6652
rect 11356 -7178 14084 -6708
<< metal5 >>
rect -2060 -6624 1008 -6518
rect -5599 -6652 1008 -6624
rect -5599 -7070 -1906 -6652
rect 796 -7070 1008 -6652
rect -5599 -7208 1008 -7070
rect 11210 -6629 14266 -6598
rect 11210 -6708 17133 -6629
rect 11210 -7178 11356 -6708
rect 14084 -7178 17133 -6708
rect 11210 -7207 17133 -7178
rect -5599 -7216 -1600 -7208
rect -5599 -9230 -5007 -7216
rect 11210 -7274 14266 -7207
rect 16555 -9228 17133 -7207
rect -5599 -9232 -4904 -9230
rect -5599 -9236 -3578 -9232
rect -5600 -9238 -3578 -9236
rect -5600 -9812 -3414 -9238
rect 3356 -9804 8142 -9236
rect 15434 -9806 17133 -9228
rect -5600 -9820 -3578 -9812
rect -5599 -9822 -3578 -9820
rect -5599 -9828 -4218 -9822
rect -5599 -11320 -5025 -9828
rect 16555 -11312 17133 -9806
rect -5599 -11904 -3670 -11320
rect 3372 -11894 8158 -11326
rect 15396 -11892 17133 -11312
rect -5599 -13422 -5025 -11904
rect 16555 -13392 17133 -11892
rect -4350 -13422 -3458 -13396
rect -5606 -13978 -3458 -13422
rect 3232 -13978 8170 -13398
rect 15374 -13972 17133 -13392
rect -5599 -15516 -5025 -13978
rect -4350 -13980 -3458 -13978
rect 16555 -15482 17133 -13972
rect -5610 -16072 -3680 -15516
rect 3378 -16066 8316 -15486
rect 15308 -16062 17133 -15482
rect -5599 -17588 -5025 -16072
rect 16555 -17564 17133 -16062
rect -5599 -18144 -3624 -17588
rect 3328 -18144 8266 -17564
rect 15326 -18144 17133 -17564
rect -5599 -19678 -5025 -18144
rect -5599 -20232 -3434 -19678
rect 3372 -20224 8310 -19644
rect 16555 -19646 17133 -18144
rect 15294 -20226 17133 -19646
rect -5599 -20234 -3614 -20232
rect -5599 -21762 -5025 -20234
rect 16555 -21735 17133 -20226
rect -5599 -22318 -3432 -21762
rect -5599 -23834 -5025 -22318
rect 3384 -22324 8322 -21744
rect 15297 -22313 17133 -21735
rect -5599 -24404 -3418 -23834
rect -5599 -24408 -3632 -24404
rect 3396 -24408 8334 -23828
rect 16555 -23839 17133 -22313
rect -5599 -29031 -5025 -24408
rect 15223 -24417 17133 -23839
rect -5599 -29605 4737 -29031
use capacitors_5  capacitors_5_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698317566
transform 1 0 -3998 0 1 -9812
box -32 -14934 9494 2050
use capacitors_5  capacitors_5_1
timestamp 1698317566
transform -1 0 15592 0 1 -9806
box -32 -14934 9494 2050
use clock  clock_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698240185
transform 0 -1 5624 1 0 -32914
box -410 -1832 6030 1274
use nmos_diode2  nmos_diode2_0
timestamp 1698329102
transform 1 0 4962 0 1 -24914
box -46 -1200 1674 106
use nmos_dnw2  nmos_dnw2_0
timestamp 1698328972
transform 1 0 5430 0 1 -8420
box -466 818 1510 2262
<< labels >>
rlabel space 5400 -7370 5400 -7370 1 vin
rlabel metal1 5360 -7478 5360 -7478 1 vin
port 1 n
rlabel metal1 4550 -7416 4550 -7416 1 vs
port 2 n
rlabel metal3 5666 -7662 5666 -7662 1 node1
port 3 n
rlabel metal3 5980 -7712 5980 -7712 1 node2
port 4 n
rlabel metal2 5176 -8760 5176 -8760 1 in1
port 5 n
rlabel metal2 5624 -10848 5624 -10848 1 in2
port 6 n
rlabel metal2 5718 -12926 5718 -12926 1 in3
port 7 n
rlabel metal2 5724 -15012 5724 -15012 1 in4
port 8 n
rlabel metal2 5762 -17098 5762 -17098 1 in5
port 9 n
rlabel metal2 5660 -19180 5660 -19180 1 in6
port 10 n
rlabel metal2 5798 -21270 5798 -21270 1 in7
port 11 n
rlabel metal2 5728 -23350 5728 -23350 1 in8
port 12 n
rlabel metal1 5762 -25952 5762 -25952 1 out
port 13 n
rlabel metal1 5578 -26838 5578 -26838 1 clk
port 14 n
rlabel metal1 5934 -26832 5934 -26832 1 clkb
port 15 n
rlabel metal5 3780 -29232 3780 -29232 1 gnd
port 16 n
rlabel metal4 8228 -28904 8228 -28904 1 vdd
port 17 n
rlabel metal1 3328 -11112 3328 -11112 1 clk_in1
port 18 n
rlabel metal1 3374 -23414 3374 -23414 1 clk_in3
port 20 n
rlabel poly 5526 -6336 5526 -6336 1 gate1
rlabel poly 6116 -6348 6116 -6348 1 gate2
<< end >>
