magic
tech sky130A
magscale 1 2
timestamp 1697813608
<< locali >>
rect 2418 3684 4121 3693
rect 2418 3646 3518 3647
rect 2418 3625 2604 3646
rect 2672 3516 2742 3644
rect 2876 3625 3518 3646
rect 3598 3625 4121 3647
rect 3836 3520 3900 3625
rect 2806 3434 2890 3436
rect 3658 3434 3964 3440
rect 2806 3433 3034 3434
rect 2634 3392 3034 3433
rect 3544 3392 3964 3434
rect 3658 3385 3964 3392
rect 3658 3384 3730 3385
rect 1774 3248 1868 3384
rect 3894 3382 3964 3385
rect 2224 2970 2318 3106
rect 4256 2970 4350 3106
rect 2474 2916 2624 2922
rect 1900 2836 2050 2900
rect 2474 2858 2738 2916
rect 3960 2906 4080 2912
rect 3960 2902 4090 2906
rect 3852 2854 4090 2902
rect 3852 2844 4080 2854
rect 3960 2840 4080 2844
rect 4524 2840 4678 2924
rect 2420 2690 2938 2692
rect 3054 2690 4123 2692
rect 2420 2672 4123 2690
rect 4122 2635 4123 2672
rect 2420 2624 4123 2635
<< viali >>
rect 2415 3650 4123 3684
rect 2415 3647 3518 3650
rect 3598 3647 4123 3650
rect 2414 2635 4122 2672
<< metal1 >>
rect 2418 3690 4121 3693
rect 2403 3684 4135 3690
rect 2403 3647 2415 3684
rect 3518 3647 3598 3650
rect 4123 3647 4135 3684
rect 2403 3641 4135 3647
rect 2418 3626 4121 3641
rect 2418 3625 3518 3626
rect 3598 3625 4121 3626
rect 2598 3624 2916 3625
rect 2971 3624 3010 3625
rect 3737 3622 3775 3625
rect 3146 3374 3250 3432
rect 3212 2934 3250 3374
rect 3182 2919 3250 2934
rect 3148 2918 3250 2919
rect 3136 2832 3146 2918
rect 3204 2844 3250 2918
rect 3307 3393 3410 3432
rect 3307 2897 3346 3393
rect 3307 2844 3319 2897
rect 3204 2832 3222 2844
rect 3148 2830 3222 2832
rect 3309 2830 3319 2844
rect 3392 2883 3402 2897
rect 3392 2844 3414 2883
rect 3392 2830 3402 2844
rect 3062 2760 3510 2797
rect 1412 2618 1422 2700
rect 1496 2618 1506 2700
rect 2678 2693 2713 2696
rect 2418 2690 2938 2693
rect 3054 2692 3510 2693
rect 3958 2692 4121 2693
rect 3054 2690 4121 2692
rect 2418 2678 4121 2690
rect 1818 2672 4134 2678
rect 1818 2635 2414 2672
rect 4122 2635 4134 2672
rect 1818 2629 4134 2635
rect 2418 2625 4121 2629
rect 5504 2372 5514 2448
rect 5598 2372 5608 2448
<< via1 >>
rect 3146 2832 3204 2918
rect 3319 2830 3392 2897
rect 1422 2618 1496 2700
rect 5514 2372 5598 2448
<< metal2 >>
rect 3146 2918 3204 2928
rect 3319 2897 3392 2907
rect 3146 2822 3204 2832
rect 3307 2830 3319 2857
rect 1402 2724 1516 2734
rect 3158 2678 3198 2822
rect 1516 2638 3198 2678
rect 3307 2820 3392 2830
rect 1402 2602 1516 2612
rect 3307 2614 3348 2820
rect 3307 2573 5598 2614
rect 5557 2468 5598 2573
rect 5484 2458 5600 2468
rect 5484 2346 5600 2356
<< via2 >>
rect 1402 2700 1516 2724
rect 1402 2618 1422 2700
rect 1422 2618 1496 2700
rect 1496 2618 1516 2700
rect 1402 2612 1516 2618
rect 5484 2448 5600 2458
rect 5484 2372 5514 2448
rect 5514 2372 5598 2448
rect 5598 2372 5600 2448
rect 5484 2356 5600 2372
<< metal3 >>
rect 1376 2608 1386 2748
rect 1536 2608 1546 2748
rect 1392 2607 1526 2608
rect 5474 2458 5610 2463
rect 5474 2356 5484 2458
rect 5600 2356 5610 2458
rect 5474 2351 5610 2356
<< via3 >>
rect 1386 2724 1536 2748
rect 1386 2612 1402 2724
rect 1402 2612 1516 2724
rect 1516 2612 1536 2724
rect 1386 2608 1536 2612
<< metal4 >>
rect 1385 2748 1537 2749
rect 1385 2608 1386 2748
rect 1536 2608 1537 2748
rect 1385 2607 1537 2608
rect 1410 2226 1494 2607
use sky130_fd_pr__nfet_01v8_U3V43Z  sky130_fd_pr__nfet_01v8_U3V43Z_0
timestamp 1697813328
transform 1 0 2261 0 1 2882
box -396 -260 396 260
use sky130_fd_pr__nfet_01v8_U3V43Z  sky130_fd_pr__nfet_01v8_U3V43Z_1
timestamp 1697813328
transform 1 0 4319 0 1 2882
box -396 -260 396 260
use sky130_fd_pr__pfet_01v8_lvt_TM5SY6  sky130_fd_pr__pfet_01v8_lvt_TM5SY6_0
timestamp 1697811387
transform 1 0 3868 0 1 3424
box -246 -269 246 269
use sky130_fd_pr__cap_mim_m3_1_TNHPNJ  XC3
timestamp 1697379271
transform 1 0 3433 0 1 1481
box -2186 -1040 2186 1040
use sky130_fd_pr__nfet_01v8_U3V43Z  XM1
timestamp 1697813328
transform 1 0 2947 0 1 2882
box -396 -260 396 260
use sky130_fd_pr__nfet_01v8_U3V43Z  XM2
timestamp 1697813328
transform 1 0 3633 0 1 2882
box -396 -260 396 260
use sky130_fd_pr__pfet_01v8_lvt_TM5SY6  XM3
timestamp 1697811387
transform 1 0 3482 0 1 3424
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_lvt_TM5SY6  XM6
timestamp 1697811387
transform 1 0 2710 0 1 3424
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_lvt_TM5SY6  XM18
timestamp 1697811387
transform 1 0 3096 0 1 3424
box -246 -269 246 269
<< labels >>
rlabel metal2 4602 2614 4602 2614 1 vo1
rlabel metal1 4056 3693 4056 3693 1 Vdd
rlabel metal1 4134 2653 4134 2653 3 gnd
<< end >>
