magic
tech sky130A
magscale 1 2
timestamp 1698622305
<< nwell >>
rect -246 -269 246 269
<< pmoslvt >>
rect -50 -50 50 50
<< pdiff >>
rect -108 38 -50 50
rect -108 -38 -96 38
rect -62 -38 -50 38
rect -108 -50 -50 -38
rect 50 38 108 50
rect 50 -38 62 38
rect 96 -38 108 38
rect 50 -50 108 -38
<< pdiffc >>
rect -96 -38 -62 38
rect 62 -38 96 38
<< nsubdiff >>
rect -210 199 -114 233
rect 114 199 210 233
rect -210 137 -176 199
rect 176 137 210 199
rect -210 -199 -176 -137
rect 176 -199 210 -137
rect -210 -233 -114 -199
rect 114 -233 210 -199
<< nsubdiffcont >>
rect -114 199 114 233
rect -210 -137 -176 137
rect 176 -137 210 137
rect -114 -233 114 -199
<< poly >>
rect -50 131 50 147
rect -50 97 -34 131
rect 34 97 50 131
rect -50 50 50 97
rect -50 -97 50 -50
rect -50 -131 -34 -97
rect 34 -131 50 -97
rect -50 -147 50 -131
<< polycont >>
rect -34 97 34 131
rect -34 -131 34 -97
<< locali >>
rect -210 199 -114 233
rect 114 199 210 233
rect -210 137 -176 199
rect 176 137 210 199
rect -50 97 -34 131
rect 34 97 50 131
rect -96 38 -62 54
rect -96 -54 -62 -38
rect 62 38 96 54
rect 62 -54 96 -38
rect -50 -131 -34 -97
rect 34 -131 50 -97
rect -210 -199 -176 -137
rect 176 -199 210 -137
rect -210 -233 -114 -199
rect 114 -233 210 -199
<< viali >>
rect -34 97 34 131
rect -96 -38 -62 38
rect 62 -38 96 38
rect -34 -131 34 -97
<< metal1 >>
rect -46 131 46 137
rect -46 97 -34 131
rect 34 97 46 131
rect -46 91 46 97
rect -102 38 -56 50
rect -102 -38 -96 38
rect -62 -38 -56 38
rect -102 -50 -56 -38
rect 56 38 102 50
rect 56 -38 62 38
rect 96 -38 102 38
rect 56 -50 102 -38
rect -46 -97 46 -91
rect -46 -131 -34 -97
rect 34 -131 46 -97
rect -46 -137 46 -131
<< properties >>
string FIXED_BBOX -193 -216 193 216
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
