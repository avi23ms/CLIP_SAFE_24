magic
tech sky130A
magscale 1 2
timestamp 1698416676
<< error_s >>
rect 2722 488 2755 524
rect 2756 522 2789 524
rect 1192 414 1314 435
rect 1580 418 1700 435
rect 1194 386 1286 407
rect 1580 390 1672 407
rect 2720 -2026 2753 -1990
rect 2754 -1992 2787 -1990
rect 1190 -2100 1312 -2079
rect 1578 -2096 1698 -2079
rect 1192 -2128 1284 -2107
rect 1578 -2124 1670 -2107
<< metal1 >>
rect -4 2064 6228 2128
rect -22 1860 -12 2064
rect 6214 1860 6228 2064
rect -4 1774 6228 1860
rect 5723 1687 5843 1774
rect 5960 1747 6076 1774
rect 5724 641 5840 1687
rect 5251 499 5842 641
rect 5724 -1866 5840 499
rect 5338 -1985 5840 -1866
rect 5338 -2003 5839 -1985
rect 5366 -3170 5520 -3166
rect -16 -3274 5742 -3170
rect -16 -3344 6206 -3274
rect 8 -3390 6206 -3344
rect 0 -3568 10 -3390
rect 6176 -3568 6206 -3390
rect 8 -3668 6206 -3568
<< via1 >>
rect -12 1860 6214 2064
rect 10 -3568 6176 -3390
<< metal2 >>
rect -12 2064 6214 2074
rect -12 1850 6214 1860
rect 10 -3390 6176 -3380
rect 10 -3578 6176 -3568
<< via2 >>
rect -12 1860 6214 2064
rect 10 -3568 6176 -3390
<< metal3 >>
rect -22 1824 -12 2106
rect 6220 1824 6230 2106
rect 0 -3568 10 -3350
rect 6172 -3385 6182 -3350
rect 6172 -3390 6186 -3385
rect 6176 -3568 6186 -3390
rect 0 -3573 6186 -3568
<< via3 >>
rect -12 2064 6220 2106
rect -12 1860 6214 2064
rect 6214 1860 6220 2064
rect -12 1824 6220 1860
rect 10 -3390 6172 -3350
rect 10 -3568 6172 -3390
<< metal4 >>
rect -12 2107 6242 2144
rect -13 2106 6242 2107
rect -13 1824 -12 2106
rect 6220 1824 6242 2106
rect -13 1823 6242 1824
rect -12 1747 6242 1823
rect -12 1744 5229 1747
rect 5885 1744 6242 1747
rect 9 -3350 26 -3349
rect 9 -3568 10 -3350
rect 9 -3569 26 -3568
<< via4 >>
rect 26 -3350 6178 -3346
rect 26 -3568 6172 -3350
rect 6172 -3568 6178 -3350
rect 26 -3628 6178 -3568
<< metal5 >>
rect 8 -3322 6204 -3268
rect 2 -3346 6204 -3322
rect 2 -3628 26 -3346
rect 6178 -3628 6204 -3346
rect 2 -3652 6204 -3628
rect 8 -3668 6204 -3652
use comparator_full  comparator_full_0
timestamp 1698416676
transform 1 0 166 0 1 -756
box -8 -5 5299 2483
use comparator_full  comparator_full_1
timestamp 1698416676
transform 1 0 164 0 1 -3270
box -8 -5 5299 2483
<< end >>
