magic
tech sky130A
magscale 1 2
timestamp 1698771642
<< nwell >>
rect -494 -164 494 198
<< pmoslvt >>
rect -400 -64 400 136
<< pdiff >>
rect -458 124 -400 136
rect -458 -52 -446 124
rect -412 -52 -400 124
rect -458 -64 -400 -52
rect 400 124 458 136
rect 400 -52 412 124
rect 446 -52 458 124
rect 400 -64 458 -52
<< pdiffc >>
rect -446 -52 -412 124
rect 412 -52 446 124
<< poly >>
rect -400 136 400 162
rect -400 -111 400 -64
rect -400 -145 -384 -111
rect 384 -145 400 -111
rect -400 -161 400 -145
<< polycont >>
rect -384 -145 384 -111
<< locali >>
rect -446 124 -412 140
rect -446 -68 -412 -52
rect 412 124 446 140
rect 412 -68 446 -52
rect -400 -145 -384 -111
rect 384 -145 400 -111
<< viali >>
rect -446 -52 -412 124
rect 412 -52 446 124
rect -384 -145 384 -111
<< metal1 >>
rect -452 124 -406 136
rect -452 -52 -446 124
rect -412 -52 -406 124
rect -452 -64 -406 -52
rect 406 124 452 136
rect 406 -52 412 124
rect 446 -52 452 124
rect 406 -64 452 -52
rect -396 -111 396 -105
rect -396 -145 -384 -111
rect 384 -145 396 -111
rect -396 -151 396 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 4 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
