magic
tech sky130A
magscale 1 2
timestamp 1698416676
<< error_s >>
rect 2556 1244 2589 1280
rect 2590 1278 2623 1280
rect 1026 1170 1148 1191
rect 1414 1174 1534 1191
rect 1028 1142 1120 1163
rect 1414 1146 1506 1163
<< locali >>
rect 890 1654 916 2275
rect 958 2046 974 2275
rect 958 1990 986 2046
rect 958 1654 974 1990
rect 890 1638 974 1654
rect 2558 1382 2914 1384
rect 824 1312 894 1382
rect 2558 1280 2946 1382
rect 2590 1278 2946 1280
rect 2778 -3 2905 107
<< viali >>
rect 1695 2411 2052 2448
rect 916 1654 958 2275
<< metal1 >>
rect 40 2470 2056 2471
rect -8 2464 2056 2470
rect -8 2448 2063 2464
rect -8 2423 1695 2448
rect -8 -5 40 2423
rect 1687 2411 1695 2423
rect 2052 2411 2063 2448
rect 1687 2398 2063 2411
rect 888 2275 975 2287
rect 888 2194 916 2275
rect 890 1706 916 2194
rect 886 1654 916 1706
rect 958 2194 975 2275
rect 958 1706 974 2194
rect 1374 2190 1384 2296
rect 1438 2190 1448 2296
rect 2009 2267 4931 2270
rect 2009 2209 4220 2267
rect 4821 2209 4931 2267
rect 2009 2200 4931 2209
rect 2139 2164 3290 2166
rect 2135 2162 3290 2164
rect 1130 2148 3290 2162
rect 1130 2098 2779 2148
rect 2135 2094 2779 2098
rect 3272 2094 3290 2148
rect 2135 2071 3290 2094
rect 3105 2070 3290 2071
rect 2060 1904 3038 1908
rect 2060 1902 2594 1904
rect 1002 1816 1012 1882
rect 1100 1816 1110 1882
rect 2012 1824 2594 1902
rect 3029 1824 3039 1904
rect 2012 1814 3038 1824
rect 4026 1772 4036 1780
rect 958 1654 978 1706
rect 1130 1689 4036 1772
rect 4536 1689 4546 1780
rect 1130 1686 4540 1689
rect 886 1386 978 1654
rect 226 1270 3190 1386
rect 3340 1270 3609 1386
rect 3723 1270 4616 1386
rect 4860 1270 5109 1386
rect 1026 1170 1036 1236
rect 1140 1170 1150 1236
rect 1414 1174 1424 1238
rect 1524 1174 1534 1238
rect 4484 1163 4494 1240
rect 4610 1163 4620 1240
rect 4122 652 4170 686
rect 196 478 284 512
rect 592 476 680 510
rect 1762 478 1850 512
rect 2142 478 2230 512
rect 950 364 960 428
rect 1020 364 1030 428
rect 1330 352 1340 412
rect 1396 352 1406 412
rect 1718 356 1728 410
rect 1786 356 1796 410
rect 2098 364 2108 420
rect 2160 364 2170 420
rect 1522 238 1532 292
rect 1590 238 1600 292
rect 2778 -3 2905 107
<< via1 >>
rect 1384 2190 1438 2296
rect 4220 2209 4821 2267
rect 2779 2094 3272 2148
rect 1012 1816 1100 1882
rect 2594 1824 3029 1904
rect 4036 1689 4536 1780
rect 1036 1170 1140 1236
rect 1424 1174 1524 1238
rect 4494 1163 4610 1240
rect 960 364 1020 428
rect 1340 352 1396 412
rect 1728 356 1786 410
rect 2108 364 2160 420
rect 1532 238 1590 292
<< metal2 >>
rect 1384 2296 1438 2306
rect 2051 2267 4990 2277
rect 1438 2190 1480 2256
rect 2051 2209 4220 2267
rect 4821 2209 4990 2267
rect 2051 2195 4990 2209
rect 1384 2180 1480 2190
rect 1012 1890 1100 1892
rect 1012 1882 1106 1890
rect 1100 1816 1106 1882
rect 1012 1806 1106 1816
rect 1042 1432 1106 1806
rect 1042 1246 1110 1432
rect 1436 1248 1480 2180
rect 2136 2164 3423 2166
rect 2135 2148 3423 2164
rect 2135 2094 2779 2148
rect 3272 2094 3423 2148
rect 2135 2071 3423 2094
rect 3105 2070 3290 2071
rect 2049 1904 3048 1916
rect 2049 1824 2594 1904
rect 3029 1824 3048 1904
rect 2049 1813 3048 1824
rect 1036 1236 1140 1246
rect 1036 1160 1140 1170
rect 1424 1238 1524 1248
rect 1424 1164 1524 1174
rect 2945 1161 3048 1813
rect 3327 1152 3422 2071
rect 4501 1790 4595 1796
rect 4036 1780 4595 1790
rect 4536 1689 4595 1780
rect 4036 1679 4595 1689
rect 4501 1250 4595 1679
rect 4494 1240 4610 1250
rect 4908 1173 4990 2195
rect 4494 1153 4610 1163
rect 960 428 1020 438
rect 960 354 1020 364
rect 1330 412 1400 424
rect 1730 420 1786 434
rect 1330 352 1340 412
rect 1396 352 1400 412
rect 1728 410 1786 420
rect 1330 238 1400 352
rect 1522 292 1598 402
rect 1728 346 1786 356
rect 1522 238 1532 292
rect 1590 238 1598 292
rect 1730 248 1786 346
rect 2098 420 2180 442
rect 2098 364 2108 420
rect 2160 364 2180 420
rect 2098 246 2180 364
rect 1522 234 1598 238
rect 1532 228 1590 234
use comparator_layout  comparator_layout_0
timestamp 1698405169
transform 1 0 -679 0 1 -1004
box 679 1001 3544 2340
use inverter  inverter_0
timestamp 1698167777
transform 0 -1 2178 -1 0 2429
box -54 -5 439 1260
use inverter  inverter_1
timestamp 1698167777
transform 0 -1 2178 -1 0 2043
box -54 -5 439 1260
use latch_layout  latch_layout_0
timestamp 1698416676
transform 1 0 2625 0 1 -844
box 30 840 2674 2181
<< end >>
