magic
tech sky130A
magscale 1 2
timestamp 1727000951
<< error_p >>
rect 30370 33062 30414 33098
rect 30356 33024 30394 33060
rect 58759 2350 58781 2546
rect 58819 2290 58841 2546
rect 46377 500 46465 552
rect 46411 466 46499 498
rect 70061 442 70105 456
rect 70073 404 70109 418
rect 91191 394 91279 414
rect 91189 368 91279 394
rect 91219 334 91311 360
rect 46058 71 46059 78
rect 46093 71 46277 78
rect 46311 71 46475 78
rect 49058 57 49059 78
rect 49093 57 49277 78
rect 46030 43 46059 50
rect 46093 43 46277 50
rect 46311 43 46503 50
rect 49030 29 49059 50
rect 49093 29 49277 50
rect 59963 -31521 59985 -31265
rect 60023 -31461 60045 -31265
rect 21729 -33312 21779 -33307
rect 72339 -33311 72427 -33259
rect 21757 -33340 21779 -33335
rect 72305 -33345 72393 -33313
rect 48699 -33369 48743 -33355
rect 95309 -33373 95353 -33369
rect 27525 -33417 27613 -33397
rect 48695 -33407 48731 -33393
rect 95275 -33411 95317 -33407
rect 27525 -33443 27615 -33417
rect 27493 -33477 27585 -33451
rect 69527 -33754 69711 -33733
rect 69745 -33754 69746 -33733
rect 72329 -33740 72493 -33733
rect 72527 -33740 72711 -33733
rect 72745 -33740 72746 -33733
rect 69527 -33782 69711 -33761
rect 69745 -33782 69774 -33761
rect 72301 -33768 72493 -33761
rect 72527 -33768 72711 -33761
rect 72745 -33768 72774 -33761
<< error_s >>
rect 97025 499 97075 504
rect 97025 471 97047 476
rect 23451 438 23495 442
rect 23487 400 23529 404
<< metal1 >>
rect -3290 58692 -3124 58760
rect -3290 57994 -3238 58692
rect -3154 57994 -3124 58692
rect -3610 28804 -3444 28855
rect -3634 26074 -3468 26308
rect -3634 25204 -3596 26074
rect -3502 25204 -3468 26074
rect -3634 -21452 -3468 25204
rect -3290 12352 -3124 57994
rect -2970 56598 -2822 56688
rect -2970 55900 -2936 56598
rect -2852 55900 -2822 56598
rect -2970 24162 -2822 55900
rect -2330 54500 -2164 54543
rect -2330 53802 -2294 54500
rect -2210 53802 -2164 54500
rect -2970 14472 -2804 24162
rect -2970 13612 -2946 14472
rect -2852 13612 -2804 14472
rect -2970 13483 -2804 13612
rect -2650 24058 -2484 24162
rect -2650 23188 -2606 24058
rect -2512 23188 -2484 24058
rect -3290 11492 -3238 12352
rect -3144 11492 -3124 12352
rect -3290 11482 -3124 11492
rect -2650 -19328 -2484 23188
rect -2330 16540 -2164 53802
rect -1690 52400 -1524 52474
rect -1690 51702 -1638 52400
rect -1554 51702 -1524 52400
rect -2330 15680 -2284 16540
rect -2190 15680 -2164 16540
rect -2330 15647 -2164 15680
rect -2010 21994 -1844 22016
rect -2010 21124 -1976 21994
rect -1882 21124 -1844 21994
rect -2010 -17302 -1844 21124
rect -1690 18604 -1524 51702
rect -1050 50300 -884 50353
rect -1050 49602 -1002 50300
rect -918 49602 -884 50300
rect -1050 20688 -884 49602
rect -730 48222 -564 48247
rect -730 47524 -696 48222
rect -612 47524 -564 48222
rect -730 22740 -564 47524
rect -410 46134 -244 46178
rect -410 45436 -362 46134
rect -278 45436 -244 46134
rect -410 24828 -244 45436
rect -50 44034 116 44096
rect -50 43336 2 44034
rect 86 43336 116 44034
rect -50 26906 116 43336
rect 93902 39872 95162 40182
rect 93902 39792 94104 39872
rect 93882 38954 94104 39792
rect 94960 38954 95162 39872
rect 93882 38768 95162 38954
rect 46860 29878 46996 29882
rect 46856 29814 48190 29878
rect 46856 29632 46904 29814
rect 48118 29632 48190 29814
rect 46856 29592 48190 29632
rect 46860 27902 46996 29592
rect 93336 28918 93500 28934
rect 93332 28878 93510 28918
rect 93332 28074 93374 28878
rect 93460 28074 93510 28878
rect 93332 28040 93510 28074
rect 93340 27912 93476 28040
rect 93882 27152 94010 38768
rect -50 26140 -8 26906
rect 86 26140 116 26906
rect -50 26070 116 26140
rect -410 24062 -372 24828
rect -278 24062 -244 24828
rect -410 23982 -244 24062
rect -730 21974 -684 22740
rect -590 21974 -564 22740
rect -730 21933 -564 21974
rect -1050 19922 -1018 20688
rect -924 19922 -884 20688
rect -1690 17744 -1658 18604
rect -1564 17744 -1524 18604
rect -1690 17731 -1524 17744
rect -1370 19832 -1204 19882
rect -1370 18962 -1330 19832
rect -1236 18962 -1204 19832
rect -1050 19817 -884 19922
rect -1370 -15204 -1204 18962
rect -1050 17790 -884 17808
rect -1050 16920 -1018 17790
rect -924 16920 -884 17790
rect -1050 -13132 -884 16920
rect -730 15682 -564 15704
rect -730 14812 -696 15682
rect -602 14812 -564 15682
rect -730 -11094 -564 14812
rect -410 13618 -244 13630
rect -410 12748 -368 13618
rect -274 12748 -244 13618
rect 58552 13524 58602 23889
rect -410 -7786 -244 12748
rect -50 11504 116 11542
rect -50 10634 -8 11504
rect 86 10634 116 11504
rect -50 -6878 116 10634
rect 23530 10128 24048 10240
rect 23530 9647 23594 10128
rect 22653 9576 23594 9647
rect 23942 9576 24048 10128
rect 70527 10236 70657 10243
rect 70527 10168 70712 10236
rect 70527 9655 70566 10168
rect 22653 9520 24048 9576
rect 68939 9574 70566 9655
rect 70680 9574 70712 10168
rect 68939 9530 70712 9574
rect 68939 9525 70691 9530
rect 22653 9517 23765 9520
rect 3294 -3158 4642 -3144
rect 3294 -3218 25199 -3158
rect 3294 -3414 3368 -3218
rect 4494 -3294 25199 -3218
rect 4494 -3414 4642 -3294
rect 3294 -3448 4642 -3414
rect 23874 -3794 24074 -3716
rect 23874 -4352 23912 -3794
rect 24026 -4352 24074 -3794
rect 23874 -4378 24074 -4352
rect 23938 -6659 24066 -4378
rect 25063 -5899 25199 -3294
rect 71522 -5909 71872 -5773
rect 71522 -6276 71658 -5909
rect 71430 -6318 71658 -6276
rect 71430 -6538 71468 -6318
rect 71624 -6538 71658 -6318
rect 71430 -6576 71658 -6538
rect 71522 -6580 71658 -6576
rect -50 -7722 -32 -6878
rect 82 -7722 116 -6878
rect -50 -7786 116 -7722
rect -410 -8918 -248 -7786
rect -410 -9762 -374 -8918
rect -260 -9208 -248 -8918
rect -260 -9762 -244 -9208
rect -410 -9908 -244 -9762
rect -730 -11938 -700 -11094
rect -586 -11938 -564 -11094
rect -730 -11960 -564 -11938
rect -1050 -13976 -1024 -13132
rect -910 -13976 -884 -13132
rect -1050 -14012 -884 -13976
rect -1370 -16048 -1334 -15204
rect -1220 -16048 -1204 -15204
rect -1370 -16092 -1204 -16048
rect -2010 -18146 -1980 -17302
rect -1866 -18146 -1844 -17302
rect -2010 -18224 -1844 -18146
rect -2650 -20172 -2632 -19328
rect -2518 -20172 -2484 -19328
rect -2650 -20388 -2484 -20172
rect -3634 -22296 -3614 -21452
rect -3500 -22296 -3468 -21452
rect -3634 -22438 -3468 -22296
rect 48407 -23578 48537 -23565
rect 48262 -23654 48660 -23578
rect 95011 -23604 95141 -23589
rect 48262 -24006 48300 -23654
rect 48614 -24006 48660 -23654
rect 48262 -24060 48660 -24006
rect 94916 -23698 95418 -23604
rect 48407 -24156 48537 -24060
rect 48407 -24286 49631 -24156
rect 94916 -24260 95026 -23698
rect 95340 -24164 95418 -23698
rect 95340 -24260 96615 -24164
rect 94916 -24276 96615 -24260
rect 94940 -24294 96615 -24276
rect 94940 -24328 95418 -24294
<< via1 >>
rect -3238 57994 -3154 58692
rect -3596 25204 -3502 26074
rect -2936 55900 -2852 56598
rect -2294 53802 -2210 54500
rect -2946 13612 -2852 14472
rect -2606 23188 -2512 24058
rect -3238 11492 -3144 12352
rect -1638 51702 -1554 52400
rect -2284 15680 -2190 16540
rect -1976 21124 -1882 21994
rect -1002 49602 -918 50300
rect -696 47524 -612 48222
rect -362 45436 -278 46134
rect 2 43336 86 44034
rect 94104 38954 94960 39872
rect 46904 29632 48118 29814
rect 93374 28074 93460 28878
rect -8 26140 86 26906
rect -372 24062 -278 24828
rect -684 21974 -590 22740
rect -1018 19922 -924 20688
rect -1658 17744 -1564 18604
rect -1330 18962 -1236 19832
rect -1018 16920 -924 17790
rect -696 14812 -602 15682
rect -368 12748 -274 13618
rect -8 10634 86 11504
rect 23594 9576 23942 10128
rect 70566 9574 70680 10168
rect 3368 -3414 4494 -3218
rect 23912 -4352 24026 -3794
rect 71468 -6538 71624 -6318
rect -32 -7722 82 -6878
rect -374 -9762 -260 -8918
rect -700 -11938 -586 -11094
rect -1024 -13976 -910 -13132
rect -1334 -16048 -1220 -15204
rect -1980 -18146 -1866 -17302
rect -2632 -20172 -2518 -19328
rect -3614 -22296 -3500 -21452
rect 48300 -24006 48614 -23654
rect 95026 -24260 95340 -23698
<< metal2 >>
rect -3278 58738 -3110 58754
rect -3299 58692 2097 58738
rect -3278 57994 -3238 58692
rect -3154 57994 -3110 58692
rect -3278 57922 -3110 57994
rect -2976 56632 -2808 56664
rect -2976 56598 2023 56632
rect -2976 55900 -2936 56598
rect -2852 56586 2023 56598
rect -2852 55900 -2808 56586
rect -2976 55832 -2808 55900
rect -2342 54538 -2174 54550
rect -3201 54500 4423 54538
rect -3201 54492 -2294 54500
rect -2342 53802 -2294 54492
rect -2210 54492 4423 54500
rect -2210 53802 -2174 54492
rect -2342 53718 -2174 53802
rect -1670 52444 -1502 52482
rect -1679 52400 2061 52444
rect -1679 52398 -1638 52400
rect -1670 51702 -1638 52398
rect -1554 52398 2061 52400
rect -1554 51702 -1502 52398
rect -1670 51650 -1502 51702
rect -1060 50350 -892 50368
rect -1060 50304 2087 50350
rect -1060 50300 -892 50304
rect -1060 49602 -1002 50300
rect -918 49602 -892 50300
rect -1060 49536 -892 49602
rect -732 48256 -564 48278
rect -733 48222 2071 48256
rect -733 48210 -696 48222
rect -732 47524 -696 48210
rect -612 48210 2071 48222
rect -612 47524 -564 48210
rect -732 47446 -564 47524
rect -408 46162 -240 46184
rect -408 46134 2111 46162
rect -408 45436 -362 46134
rect -278 46116 2111 46134
rect -278 45436 -240 46116
rect -408 45352 -240 45436
rect -50 44066 118 44096
rect -53 44034 2105 44066
rect -53 44020 2 44034
rect -50 43336 2 44020
rect 86 44020 2105 44034
rect 86 43336 118 44020
rect -50 43264 118 43336
rect 95011 40182 95177 42817
rect 93902 39872 95177 40182
rect 93902 38954 94104 39872
rect 94960 39613 95177 39872
rect 94960 38954 95162 39613
rect 93902 38768 95162 38954
rect 120780 30056 120864 42280
rect 128295 42196 128734 42280
rect 93410 29972 120864 30056
rect 46986 29878 70895 29880
rect 46856 29814 70895 29878
rect 46856 29632 46904 29814
rect 48118 29640 70895 29814
rect 48118 29632 48190 29640
rect 46856 29592 48190 29632
rect 70655 27608 70895 29640
rect 93410 28934 93494 29972
rect 93336 28918 93500 28934
rect 93332 28878 93500 28918
rect 93332 28074 93374 28878
rect 93460 28074 93500 28878
rect 93332 28056 93500 28074
rect 93332 28040 93496 28056
rect 23323 27356 23563 27498
rect 70655 27490 70895 27510
rect 20702 27116 23563 27356
rect 69066 27066 70895 27490
rect 120780 27292 120864 29972
rect 116432 27228 120884 27292
rect -44 26906 122 27000
rect -44 26140 -8 26906
rect 86 26140 122 26906
rect -44 26130 122 26140
rect -6742 26082 1758 26130
rect -6742 22438 -6694 26082
rect -3634 26074 -3458 26082
rect -44 26074 122 26082
rect -3634 25204 -3596 26074
rect -3502 25204 -3458 26074
rect -3634 25146 -3458 25204
rect -404 24828 -238 24932
rect -2644 24058 -2468 24112
rect -2644 24044 -2606 24058
rect -7134 22390 -6694 22438
rect -6220 23996 -2606 24044
rect -6220 21306 -6172 23996
rect -2644 23188 -2606 23996
rect -2512 24044 -2468 24058
rect -404 24062 -372 24828
rect -278 24062 -238 24828
rect -404 24044 -238 24062
rect -2512 23996 1760 24044
rect -2512 23188 -2468 23996
rect -2644 23150 -2468 23188
rect -726 22740 -560 22848
rect -2008 21994 -1832 22040
rect -2008 21950 -1976 21994
rect -7134 21258 -6172 21306
rect -5766 21902 -1976 21950
rect -5766 20208 -5718 21902
rect -2008 21124 -1976 21902
rect -1882 21950 -1832 21994
rect -726 21974 -684 22740
rect -590 21974 -560 22740
rect -726 21950 -560 21974
rect -1882 21902 1726 21950
rect -1882 21124 -1832 21902
rect -2008 21078 -1832 21124
rect -7134 20160 -5718 20208
rect -5766 20150 -5718 20160
rect -1044 20688 -878 20764
rect -1044 19922 -1018 20688
rect -924 19922 -878 20688
rect -1382 19860 -1206 19868
rect -1044 19860 -878 19922
rect -7096 19832 1786 19860
rect -7096 19812 -1330 19832
rect -7096 19134 -7048 19812
rect -7134 19086 -7048 19134
rect -1382 18962 -1330 19812
rect -1236 19812 1786 19832
rect -1236 18962 -1206 19812
rect -1382 18906 -1206 18962
rect -1700 18604 -1534 18648
rect -7134 18076 -4354 18124
rect -4402 17762 -4354 18076
rect -1700 17762 -1658 18604
rect -4402 17744 -1658 17762
rect -1564 17762 -1534 18604
rect -1060 17790 -884 17810
rect -1060 17762 -1018 17790
rect -1564 17744 -1018 17762
rect -4402 17714 -1018 17744
rect -7134 16924 -4732 16972
rect -7134 15892 -5630 15940
rect -7134 14810 -7086 14818
rect -7134 14762 -6628 14810
rect -7134 14704 -7086 14762
rect -6676 11500 -6628 14762
rect -5678 13586 -5630 15892
rect -4780 15680 -4732 16924
rect -1060 16920 -1018 17714
rect -924 17762 -884 17790
rect -924 17714 1846 17762
rect -924 16920 -884 17714
rect -1060 16848 -884 16920
rect -2320 16540 -2154 16566
rect -2320 15680 -2284 16540
rect -2190 15680 -2154 16540
rect -742 15682 -566 15726
rect -742 15680 -696 15682
rect -4780 15632 -696 15680
rect -742 14812 -696 15632
rect -602 15680 -566 15682
rect -602 15632 1832 15680
rect -602 14812 -566 15632
rect -742 14764 -566 14812
rect -2972 13612 -2946 14472
rect -2852 13612 -2806 14472
rect -2972 13586 -2806 13612
rect -398 13618 -222 13658
rect -398 13586 -368 13618
rect -5678 13538 -368 13586
rect -398 12748 -368 13538
rect -274 13586 -222 13618
rect -274 13538 1782 13586
rect -274 12748 -222 13538
rect -398 12696 -222 12748
rect -3278 12352 -3112 12398
rect -3278 11500 -3238 12352
rect -6676 11492 -3238 11500
rect -3144 11500 -3112 12352
rect -54 11504 122 11544
rect -54 11500 -8 11504
rect -3144 11492 -8 11500
rect -6676 11452 -8 11492
rect -54 10634 -8 11452
rect 86 11500 122 11504
rect 86 11452 1844 11500
rect 86 10634 122 11452
rect -54 10582 122 10634
rect 23538 10220 24056 10232
rect 70534 10230 70712 10236
rect 23538 10128 26991 10220
rect 3294 -3144 3358 9662
rect 23538 9576 23594 10128
rect 23942 10106 26991 10128
rect 70534 10168 73615 10230
rect 23942 9576 24056 10106
rect 23538 9512 24056 9576
rect 70534 9574 70566 10168
rect 70680 10116 73615 10168
rect 70680 9574 70712 10116
rect 70534 9530 70712 9574
rect 3294 -3218 4642 -3144
rect 3294 -3414 3368 -3218
rect 4494 -3414 4642 -3218
rect 3294 -3448 4642 -3414
rect 3294 -6583 3358 -3448
rect 23893 -3716 24007 9512
rect 94000 9426 94240 10262
rect 23874 -3794 24074 -3716
rect 23874 -4352 23912 -3794
rect 24026 -4352 24074 -3794
rect 23874 -4378 24074 -4352
rect 23893 -4379 24007 -4378
rect 71430 -6318 71658 -6276
rect 47909 -6579 49482 -6339
rect 71430 -6517 71468 -6318
rect 69920 -6538 71468 -6517
rect 71624 -6517 71658 -6318
rect 95241 -6452 95481 -6318
rect 71624 -6538 71668 -6517
rect 69920 -6581 71668 -6538
rect 95241 -6692 96806 -6452
rect -64 -6878 132 -6808
rect -64 -7722 -32 -6878
rect 82 -7681 132 -6878
rect 82 -7722 3062 -7681
rect -64 -7729 3062 -7722
rect -64 -7758 132 -7729
rect -410 -8918 -214 -8880
rect -410 -9762 -374 -8918
rect -260 -9762 -214 -8918
rect -410 -9767 -214 -9762
rect -410 -9815 3046 -9767
rect -410 -9830 -214 -9815
rect -750 -11094 -554 -11020
rect -750 -11938 -700 -11094
rect -586 -11861 -554 -11094
rect -586 -11909 3030 -11861
rect -586 -11938 -554 -11909
rect -750 -11970 -554 -11938
rect -1066 -13132 -870 -13066
rect -1066 -13976 -1024 -13132
rect -910 -13951 -870 -13132
rect -910 -13976 3128 -13951
rect -1066 -13999 3128 -13976
rect -1066 -14016 -870 -13999
rect -1382 -15204 -1186 -15150
rect -1382 -16048 -1334 -15204
rect -1220 -16048 -1186 -15204
rect -1382 -16049 -1186 -16048
rect -1382 -16092 3122 -16049
rect -1382 -16100 -1186 -16092
rect -876 -16097 3122 -16092
rect -2018 -17302 -1822 -17252
rect -2018 -18146 -1980 -17302
rect -1866 -18131 -1822 -17302
rect -1866 -18146 3106 -18131
rect -2018 -18179 3106 -18146
rect -2018 -18202 -1822 -18179
rect -2668 -19328 -2472 -19294
rect -2668 -20172 -2632 -19328
rect -2518 -20172 -2472 -19328
rect -2668 -20225 -2472 -20172
rect -2668 -20244 3134 -20225
rect -2636 -20273 3134 -20244
rect -3656 -21452 -3460 -21366
rect -3656 -22296 -3614 -21452
rect -3500 -22296 -3460 -21452
rect -3656 -22311 -3460 -22296
rect -3656 -22316 3118 -22311
rect -3630 -22359 3118 -22316
rect 48262 -23581 48660 -23578
rect 45869 -23654 48660 -23581
rect 45869 -23695 48300 -23654
rect 48262 -24006 48300 -23695
rect 48614 -24006 48660 -23654
rect 92109 -23604 95253 -23591
rect 92109 -23698 95418 -23604
rect 92109 -23705 95026 -23698
rect 48262 -24060 48660 -24006
rect 94916 -24260 95026 -23705
rect 95340 -24260 95418 -23698
rect 94916 -24276 95418 -24260
rect 94940 -24328 95418 -24276
<< metal3 >>
rect -6135 32356 3619 33414
rect -6135 562 -5077 32356
rect 11390 2606 11462 2610
rect -11579 8 4823 562
rect 35426 52 35498 1524
rect -6135 -33083 -5077 8
rect -6135 -34141 6745 -33083
<< metal4 >>
rect 112630 31206 120572 31774
rect 120004 -295 120572 31206
rect 101363 -953 120781 -295
rect 120004 -34106 120572 -953
rect 102427 -34276 120572 -34106
rect 102427 -34764 120453 -34276
<< metal5 >>
rect 122034 -1549 122638 30920
rect 114551 -2207 122747 -1549
rect 122034 -35492 122638 -2207
rect 115316 -36096 122638 -35492
use CP1_5_stage  CP1_5_stage_0
timestamp 1727000951
transform 1 0 332 0 1 35216
box -1718 -4908 128204 27526
use CP2_5_stage  CP2_5_stage_0
timestamp 1727000951
transform -1 0 117527 0 1 2322
box -2079 -4599 117458 28100
use CP2_5_stage  CP2_5_stage_1
timestamp 1727000951
transform 1 0 1277 0 1 -31489
box -2079 -4599 117458 28100
<< end >>
