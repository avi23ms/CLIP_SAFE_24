magic
tech sky130A
magscale 1 2
timestamp 1698771642
<< locali >>
rect 905 2310 3268 2339
rect 905 2268 955 2310
rect 3238 2268 3268 2310
rect 905 2237 3268 2268
rect 3366 1255 3506 1316
rect 679 1071 3474 1105
rect 679 1026 722 1071
rect 679 1004 3474 1026
<< viali >>
rect 955 2268 3238 2310
rect 722 1026 3474 1071
<< metal1 >>
rect 1253 2339 1290 2340
rect 2413 2339 2450 2340
rect 905 2310 3268 2339
rect 905 2268 955 2310
rect 3238 2268 3268 2310
rect 905 2237 3268 2268
rect 1253 1897 1290 2237
rect 1321 2126 1396 2181
rect 1413 1976 1423 2038
rect 1411 1896 1421 1976
rect 1484 1958 1494 2038
rect 1482 1896 1492 1958
rect 1636 1892 1673 2237
rect 1833 2028 1872 2083
rect 1803 1948 1813 2028
rect 1874 1980 1884 2028
rect 1805 1900 1815 1948
rect 1876 1900 1886 1980
rect 1308 1776 1318 1840
rect 1416 1776 1426 1840
rect 1061 1580 1673 1616
rect 852 1342 862 1434
rect 856 1290 866 1342
rect 858 1257 868 1290
rect 929 1257 939 1434
rect 1061 1257 1097 1580
rect 1239 1385 1249 1438
rect 1237 1253 1247 1385
rect 1312 1361 1322 1438
rect 1310 1253 1320 1361
rect 1444 1258 1480 1580
rect 1637 1314 1673 1580
rect 1714 1535 1788 1840
rect 1704 1482 1714 1535
rect 1793 1482 1803 1535
rect 1833 1411 1872 1900
rect 2022 1892 2059 2237
rect 2214 2034 2253 2089
rect 2194 1906 2204 2034
rect 2265 1906 2275 2034
rect 2105 1535 2179 1838
rect 2214 1691 2253 1906
rect 2413 1897 2450 2237
rect 2488 2174 2563 2183
rect 2867 2174 2877 2183
rect 2488 2128 2877 2174
rect 2932 2128 2942 2183
rect 2576 1980 2586 2038
rect 2568 1900 2578 1980
rect 2647 1958 2657 2038
rect 2963 2020 2973 2079
rect 3031 2020 3041 2079
rect 2639 1900 2649 1958
rect 2790 1899 2800 1958
rect 2858 1899 2868 1958
rect 2470 1776 2480 1840
rect 2578 1776 2588 1840
rect 2214 1552 2254 1691
rect 2606 1610 3025 1618
rect 2606 1585 3222 1610
rect 2085 1482 2095 1535
rect 2174 1482 2184 1535
rect 1807 1346 1817 1411
rect 1872 1346 1882 1411
rect 2214 1399 2253 1552
rect 1631 1251 1641 1314
rect 1706 1251 1716 1314
rect 1833 1253 1872 1346
rect 2194 1334 2204 1399
rect 2259 1334 2269 1399
rect 2014 1251 2024 1322
rect 2082 1251 2092 1322
rect 2214 1259 2253 1334
rect 2401 1253 2411 1320
rect 2470 1253 2480 1320
rect 2606 1278 2639 1585
rect 2992 1577 3222 1585
rect 2782 1253 2792 1334
rect 2855 1253 2865 1334
rect 2992 1258 3025 1577
rect 3189 1430 3222 1577
rect 3252 1483 3262 1539
rect 3346 1483 3356 1539
rect 3165 1349 3175 1430
rect 3232 1385 3242 1430
rect 1637 1249 1673 1251
rect 3169 1245 3179 1349
rect 3236 1245 3246 1385
rect 3272 1152 3282 1208
rect 3366 1152 3376 1208
rect 3407 1105 3481 1107
rect 679 1071 3481 1105
rect 679 1026 722 1071
rect 3474 1026 3481 1071
rect 679 1004 3481 1026
rect 3407 1001 3481 1004
<< via1 >>
rect 1423 1976 1484 2038
rect 1421 1958 1484 1976
rect 1421 1896 1482 1958
rect 1813 1980 1874 2028
rect 1813 1948 1876 1980
rect 1815 1900 1876 1948
rect 1318 1776 1416 1840
rect 862 1342 929 1434
rect 866 1290 929 1342
rect 868 1257 929 1290
rect 1249 1385 1312 1438
rect 1247 1361 1312 1385
rect 1247 1253 1310 1361
rect 1714 1482 1793 1535
rect 2204 1906 2265 2034
rect 2877 2128 2932 2183
rect 2586 1980 2647 2038
rect 2578 1958 2647 1980
rect 2973 2020 3031 2079
rect 2578 1900 2639 1958
rect 2800 1899 2858 1958
rect 2480 1776 2578 1840
rect 2095 1482 2174 1535
rect 1817 1346 1872 1411
rect 1641 1251 1706 1314
rect 2204 1334 2259 1399
rect 2024 1251 2082 1322
rect 2411 1253 2470 1320
rect 2792 1253 2855 1334
rect 3262 1483 3346 1539
rect 3175 1385 3232 1430
rect 3175 1349 3236 1385
rect 3179 1245 3236 1349
rect 3282 1152 3366 1208
<< metal2 >>
rect 2830 2271 3309 2306
rect 2888 2193 2923 2271
rect 2877 2183 2932 2193
rect 2877 2118 2932 2128
rect 1425 2048 1849 2076
rect 1423 2038 1849 2048
rect 2202 2048 2626 2084
rect 2973 2079 3031 2089
rect 2202 2038 2647 2048
rect 1421 1976 1423 1986
rect 1484 2028 1874 2038
rect 1484 1958 1813 2028
rect 2202 2034 2586 2038
rect 1874 1980 1876 1990
rect 1482 1948 1813 1958
rect 1482 1900 1815 1948
rect 2202 1906 2204 2034
rect 2265 1980 2586 2034
rect 2265 1906 2578 1980
rect 2814 1968 2844 2070
rect 2968 2040 2973 2078
rect 3031 2063 3062 2078
rect 3031 2031 3126 2063
rect 3031 2020 3062 2031
rect 2973 2010 3062 2020
rect 3024 2000 3062 2010
rect 2202 1902 2578 1906
rect 1482 1896 1876 1900
rect 2204 1896 2265 1902
rect 2639 1948 2647 1958
rect 2800 1958 2858 1968
rect 1421 1894 1876 1896
rect 1421 1886 1482 1894
rect 1815 1890 1876 1894
rect 2578 1890 2639 1900
rect 2800 1889 2858 1899
rect 1318 1840 1416 1850
rect 2480 1840 2578 1850
rect 1318 1766 1416 1776
rect 1336 1748 1416 1766
rect 2468 1776 2480 1836
rect 2468 1766 2578 1776
rect 2468 1748 2544 1766
rect 1336 1708 2544 1748
rect 1336 1700 1376 1708
rect 2814 1674 2844 1889
rect 1655 1646 2844 1674
rect 862 1434 929 1444
rect 1249 1438 1312 1448
rect 862 1332 866 1342
rect 866 1280 868 1290
rect 868 1247 929 1257
rect 1244 1385 1249 1437
rect 1244 1253 1247 1385
rect 1310 1351 1312 1361
rect 1655 1324 1685 1646
rect 1727 1588 2251 1618
rect 1727 1545 1762 1588
rect 1714 1535 1793 1545
rect 2095 1535 2174 1545
rect 1714 1472 1793 1482
rect 1835 1486 2095 1516
rect 1835 1421 1865 1486
rect 2095 1472 2174 1482
rect 1817 1411 1872 1421
rect 2216 1409 2251 1588
rect 1817 1336 1872 1346
rect 2204 1399 2259 1409
rect 890 1083 921 1247
rect 1244 1243 1310 1253
rect 1641 1314 1706 1324
rect 1244 1083 1275 1243
rect 1641 1241 1706 1251
rect 2014 1322 2093 1336
rect 2204 1324 2259 1334
rect 2792 1334 2855 1344
rect 2014 1251 2024 1322
rect 2082 1251 2093 1322
rect 2014 1241 2093 1251
rect 2411 1320 2470 1330
rect 2411 1243 2470 1253
rect 2792 1243 2855 1253
rect 2036 1156 2068 1241
rect 2421 1156 2453 1243
rect 2814 1156 2846 1243
rect 3094 1156 3126 2031
rect 3274 1549 3309 2271
rect 3262 1539 3346 1549
rect 3262 1473 3346 1483
rect 3175 1430 3232 1440
rect 3232 1386 3236 1395
rect 3232 1385 3239 1386
rect 3175 1339 3179 1349
rect 3236 1245 3239 1385
rect 3179 1235 3239 1245
rect 2036 1124 3126 1156
rect 2421 1123 2453 1124
rect 3208 1083 3239 1235
rect 3274 1218 3309 1473
rect 3274 1208 3366 1218
rect 3274 1173 3282 1208
rect 3282 1142 3366 1152
rect 890 1052 3239 1083
rect 890 1050 921 1052
use sky130_fd_pr__pfet_01v8_B5E2Q5  sky130_fd_pr__pfet_01v8_B5E2Q5_0
timestamp 1698771642
transform 1 0 2911 0 1 1980
box -246 -319 246 319
use sky130_fd_pr__nfet_01v8_PVEW3M  XM25
timestamp 1698771642
transform 1 0 982 0 1 1345
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM26
timestamp 1698771642
transform 1 0 1368 0 1 1345
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM27
timestamp 1698771642
transform 1 0 1754 0 1 1345
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM28
timestamp 1698771642
transform 1 0 2140 0 1 1345
box -246 -310 246 310
use sky130_fd_pr__pfet_01v8_X3YSY6  XM29
timestamp 1698771642
transform 1 0 1367 0 1 1980
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_X3YSY6  XM30
timestamp 1698771642
transform 1 0 1753 0 1 1980
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_X3YSY6  XM31
timestamp 1698771642
transform 1 0 2139 0 1 1980
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_X3YSY6  XM32
timestamp 1698771642
transform 1 0 2525 0 1 1980
box -246 -319 246 319
use sky130_fd_pr__nfet_01v8_PVEW3M  XM33
timestamp 1698771642
transform 1 0 2526 0 1 1345
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM34
timestamp 1698771642
transform 1 0 2912 0 1 1345
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM35
timestamp 1698771642
transform 1 0 3298 0 1 1345
box -246 -310 246 310
<< end >>
