magic
tech sky130A
magscale 1 2
timestamp 1698871213
<< locali >>
rect -736 1306 272 1339
rect 2558 1334 2914 1336
rect -736 1264 -715 1306
rect 226 1264 272 1306
rect 824 1264 894 1334
rect -736 1221 272 1264
rect 2558 1232 2946 1334
rect 2590 1230 2946 1232
rect -693 68 41 101
rect -693 22 -682 68
rect 4 22 41 68
rect -693 -1 41 22
rect 2778 -3 2905 107
<< viali >>
rect -715 1264 226 1306
rect -682 22 4 68
<< metal1 >>
rect -736 1338 272 1339
rect -736 1336 838 1338
rect -736 1306 3190 1336
rect -736 1264 -715 1306
rect 226 1264 3190 1306
rect -736 1233 3190 1264
rect -736 1222 1016 1233
rect 1568 1222 3190 1233
rect 3340 1222 3609 1336
rect 3723 1222 4470 1336
rect 5047 1222 5109 1336
rect -736 1221 272 1222
rect -527 1123 -517 1182
rect -421 1123 -411 1182
rect -143 1118 -133 1185
rect -23 1179 -13 1185
rect -22 1121 -12 1179
rect -23 1118 -13 1121
rect 1024 1115 1034 1173
rect 1145 1115 1155 1173
rect 1409 1119 1419 1189
rect 1527 1119 1537 1189
rect 4486 1121 4496 1182
rect 4618 1121 4628 1182
rect -621 1054 -529 1065
rect -625 893 -615 1054
rect -554 893 -529 1054
rect -222 1053 -156 1066
rect -225 896 -215 1053
rect -162 896 -152 1053
rect -621 888 -529 893
rect -222 887 -156 896
rect 3856 762 3882 788
rect 4062 754 4072 776
rect 4122 652 4170 686
rect 196 478 284 512
rect 1762 510 1850 512
rect 592 476 680 510
rect 1750 478 1850 510
rect 2126 478 2230 512
rect 1750 476 1804 478
rect 950 364 960 428
rect 1020 364 1030 428
rect 1330 352 1340 412
rect 1396 352 1406 412
rect 1718 356 1728 410
rect 1786 356 1796 410
rect 2098 364 2108 420
rect 2160 364 2170 420
rect 1522 238 1532 292
rect 1590 238 1600 292
rect -693 74 41 101
rect -694 68 41 74
rect -694 22 -682 68
rect 4 22 41 68
rect -694 16 41 22
rect -693 -1 41 16
rect 2778 -3 2905 107
<< via1 >>
rect -517 1123 -421 1182
rect -133 1179 -23 1185
rect -133 1121 -22 1179
rect -133 1118 -23 1121
rect 1034 1115 1145 1173
rect 1419 1119 1527 1189
rect 4496 1121 4618 1182
rect -615 893 -554 1054
rect -215 896 -162 1053
rect 960 364 1020 428
rect 1340 352 1396 412
rect 1728 356 1786 410
rect 2108 364 2160 420
rect 1532 238 1590 292
<< metal2 >>
rect -794 1463 4556 1494
rect -794 835 -763 1463
rect -601 1402 3393 1433
rect -601 1065 -570 1402
rect 1043 1336 3041 1366
rect 3362 1336 3393 1402
rect 1043 1330 3048 1336
rect -512 1201 -402 1211
rect -517 1182 -512 1192
rect -517 1121 -512 1123
rect -517 1113 -402 1121
rect -512 1111 -402 1113
rect -133 1189 -23 1191
rect -133 1185 -22 1189
rect -23 1179 -22 1185
rect 1043 1183 1079 1330
rect 1418 1198 1528 1208
rect 1034 1173 1145 1183
rect -22 1121 1034 1155
rect -23 1119 1034 1121
rect -23 1118 -22 1119
rect -133 1111 -22 1118
rect -133 1108 -23 1111
rect 1034 1105 1145 1115
rect 2945 1161 3048 1330
rect 3327 1152 3422 1336
rect 4525 1192 4556 1463
rect 4496 1182 4618 1192
rect 3362 1124 3393 1152
rect 1418 1108 1528 1118
rect 4496 1111 4618 1121
rect 4887 1188 4982 1198
rect 4887 1110 4982 1120
rect -621 1054 -529 1065
rect -621 893 -615 1054
rect -554 893 -529 1054
rect -222 1053 -156 1066
rect -222 930 -215 1053
rect -621 888 -529 893
rect -227 896 -215 930
rect -162 896 -156 1053
rect -615 883 -554 888
rect -227 887 -156 896
rect -227 886 -162 887
rect -227 835 -196 886
rect -794 804 -196 835
rect 2596 684 2628 848
rect 960 428 1020 438
rect 960 354 1020 364
rect 1330 412 1400 424
rect 1730 420 1786 434
rect 1330 352 1340 412
rect 1396 352 1400 412
rect 1728 410 1786 420
rect 1330 238 1400 352
rect 1522 292 1598 402
rect 1728 346 1786 356
rect 1522 238 1532 292
rect 1590 238 1598 292
rect 1730 248 1786 346
rect 2098 420 2180 442
rect 2098 364 2108 420
rect 2160 364 2180 420
rect 2098 246 2180 364
rect 1522 234 1598 238
rect 1532 228 1590 234
<< via2 >>
rect -512 1182 -402 1201
rect -512 1123 -421 1182
rect -421 1123 -402 1182
rect -512 1121 -402 1123
rect 1418 1189 1528 1198
rect 1418 1119 1419 1189
rect 1419 1119 1527 1189
rect 1527 1119 1528 1189
rect 1418 1118 1528 1119
rect 4887 1120 4982 1188
<< metal3 >>
rect -490 1262 4949 1323
rect -490 1206 -392 1262
rect -522 1201 -392 1206
rect -522 1121 -512 1201
rect -402 1121 -392 1201
rect 1342 1198 1538 1262
rect 1342 1122 1418 1198
rect -522 1116 -392 1121
rect 1408 1118 1418 1122
rect 1528 1118 1538 1198
rect 4888 1193 4949 1262
rect 1408 1113 1538 1118
rect 4877 1188 4992 1193
rect 4877 1120 4887 1188
rect 4982 1120 4992 1188
rect 4877 1115 4992 1120
use comparator_layout  comparator_layout_0
timestamp 1698771642
transform 1 0 -679 0 1 -1004
box 679 1001 3544 2340
use inverter  inverter_0
timestamp 1698871213
transform -1 0 110 0 1 36
box -54 -5 439 1260
use inverter  inverter_1
timestamp 1698871213
transform -1 0 -276 0 1 36
box -54 -5 439 1260
use latch_layout  latch_layout_0
timestamp 1698771642
transform 1 0 2625 0 1 -844
box 30 840 2674 2181
<< labels >>
rlabel metal2 929 1136 929 1136 1 vo-
rlabel metal3 1391 1179 1391 1179 1 vo+
rlabel via1 -595 953 -595 953 1 vo1+
rlabel via1 -204 935 -204 935 1 vo1-
rlabel metal1 2650 1244 2650 1244 1 Vdd
port 1 n
rlabel metal1 2844 16 2844 16 1 gnd
port 2 n
rlabel metal2 2612 750 2612 750 1 clk
port 3 n
rlabel metal1 2134 494 2134 494 1 Vc-
port 4 n
rlabel metal1 606 486 606 486 1 V+
port 5 n
rlabel metal1 1762 486 1762 486 1 V-
port 6 n
rlabel metal1 220 492 220 492 1 Vc+
port 7 n
rlabel metal1 3864 766 3864 766 1 Q
port 8 n
rlabel metal1 4064 760 4064 760 1 Q1
port 9 n
<< end >>
