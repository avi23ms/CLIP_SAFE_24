magic
tech sky130A
magscale 1 2
timestamp 1698404476
<< dnwell >>
rect -254 2142 1076 2232
rect -254 2048 1214 2142
rect -400 2042 1214 2048
rect -400 2034 1402 2042
rect -418 2032 1402 2034
rect -418 1130 1408 2032
rect -254 1128 1408 1130
rect -254 1020 1214 1128
rect -254 906 1076 1020
<< nwell >>
rect 1070 2256 1510 2262
rect -424 2040 1510 2256
rect -424 1130 -252 2040
rect 1070 2036 1510 2040
rect 1238 1134 1510 2036
rect 1046 1132 1510 1134
rect 748 1130 1510 1132
rect -424 896 1510 1130
rect -194 894 1510 896
rect 1070 886 1510 894
<< nmos >>
rect 80 1858 110 1942
rect 668 1858 698 1942
rect 0 1200 200 1800
rect 590 1200 790 1800
<< ndiff >>
rect 20 1920 80 1942
rect 20 1882 30 1920
rect 64 1882 80 1920
rect 20 1858 80 1882
rect 110 1928 172 1942
rect 110 1872 124 1928
rect 158 1872 172 1928
rect 110 1858 172 1872
rect 606 1928 668 1942
rect 606 1872 620 1928
rect 654 1872 668 1928
rect 606 1858 668 1872
rect 698 1920 758 1942
rect 698 1882 714 1920
rect 748 1882 758 1920
rect 698 1858 758 1882
rect -110 1770 0 1800
rect -110 1230 -90 1770
rect -40 1230 0 1770
rect -110 1200 0 1230
rect 200 1770 310 1800
rect 200 1230 230 1770
rect 280 1230 310 1770
rect 200 1200 310 1230
rect 480 1770 590 1800
rect 480 1230 510 1770
rect 560 1230 590 1770
rect 480 1200 590 1230
rect 790 1770 900 1800
rect 790 1230 830 1770
rect 880 1230 900 1770
rect 790 1200 900 1230
<< ndiffc >>
rect 30 1882 64 1920
rect 124 1872 158 1928
rect 620 1872 654 1928
rect 714 1882 748 1920
rect -90 1230 -40 1770
rect 230 1230 280 1770
rect 510 1230 560 1770
rect 830 1230 880 1770
<< psubdiff >>
rect 1048 1540 1174 1562
rect 1048 1216 1090 1540
rect 1128 1216 1174 1540
rect 1048 1198 1174 1216
<< nsubdiff >>
rect 1324 1512 1434 1544
rect 1324 1230 1348 1512
rect 1402 1230 1434 1512
rect 1324 1214 1434 1230
<< psubdiffcont >>
rect 1090 1216 1128 1540
<< nsubdiffcont >>
rect 1348 1230 1402 1512
<< poly >>
rect 80 1942 110 1972
rect 668 1942 698 1972
rect 80 1826 110 1858
rect 668 1826 698 1858
rect 0 1800 200 1826
rect 590 1800 790 1826
rect 0 1172 200 1200
rect 590 1174 790 1200
<< locali >>
rect 22 1936 72 1948
rect 20 1924 74 1936
rect 64 1878 74 1924
rect 20 1864 74 1878
rect 114 1928 170 1944
rect 114 1872 124 1928
rect 158 1872 170 1928
rect 22 1856 72 1864
rect 114 1854 170 1872
rect 608 1928 664 1944
rect 608 1872 620 1928
rect 654 1872 664 1928
rect 608 1854 664 1872
rect 704 1920 754 1946
rect 704 1882 714 1920
rect 748 1882 754 1920
rect 704 1854 754 1882
rect -108 1770 -2 1804
rect -108 1230 -90 1770
rect -40 1768 -2 1770
rect -38 1232 -2 1768
rect 202 1770 302 1796
rect 202 1768 230 1770
rect 202 1734 228 1768
rect -40 1230 -2 1232
rect -108 1190 -2 1230
rect 210 1234 228 1734
rect 280 1734 302 1770
rect 480 1790 578 1800
rect 480 1770 580 1790
rect 480 1766 510 1770
rect 480 1758 508 1766
rect 210 1230 230 1234
rect 280 1230 300 1734
rect 210 1210 300 1230
rect 490 1234 508 1758
rect 490 1230 510 1234
rect 560 1230 580 1770
rect 490 1210 580 1230
rect 790 1770 902 1818
rect 790 1230 830 1770
rect 880 1768 902 1770
rect 882 1232 902 1768
rect 880 1230 902 1232
rect 790 1204 902 1230
rect 1048 1560 1174 1562
rect 1048 1540 1464 1560
rect 1048 1216 1090 1540
rect 1128 1512 1464 1540
rect 1128 1230 1348 1512
rect 1402 1230 1464 1512
rect 1128 1216 1464 1230
rect 1048 1198 1464 1216
<< viali >>
rect 20 1920 64 1924
rect 20 1882 30 1920
rect 30 1882 64 1920
rect 20 1878 64 1882
rect 124 1872 158 1928
rect 620 1872 654 1928
rect 714 1882 748 1920
rect -90 1232 -40 1768
rect -40 1232 -38 1768
rect 228 1234 230 1768
rect 230 1234 280 1768
rect 508 1234 510 1766
rect 510 1234 560 1766
rect 830 1232 880 1768
rect 880 1232 882 1768
<< metal1 >>
rect 22 1936 72 1948
rect -114 1924 74 1936
rect -114 1878 20 1924
rect 64 1878 74 1924
rect -114 1864 74 1878
rect 114 1928 170 1946
rect 114 1872 124 1928
rect 158 1872 170 1928
rect -114 1786 -12 1864
rect 22 1856 72 1864
rect 114 1854 170 1872
rect 608 1928 664 1944
rect 608 1872 620 1928
rect 654 1872 664 1928
rect 608 1854 664 1872
rect 704 1936 754 1946
rect 704 1920 902 1936
rect 704 1882 714 1920
rect 748 1882 902 1920
rect 704 1864 902 1882
rect 704 1854 754 1864
rect 802 1862 902 1864
rect -114 1768 -2 1786
rect -114 1232 -90 1768
rect -38 1232 -2 1768
rect -114 1210 -2 1232
rect 200 1772 312 1802
rect 200 1230 210 1772
rect 302 1230 312 1772
rect 480 1772 590 1800
rect 802 1798 904 1862
rect 480 1269 494 1772
rect -114 1104 -12 1210
rect 200 1202 312 1230
rect 479 1230 494 1269
rect 576 1230 590 1772
rect 479 1202 590 1230
rect 794 1768 904 1798
rect 794 1232 830 1768
rect 882 1232 904 1768
rect 794 1208 904 1232
rect 210 1190 300 1202
rect 479 1190 569 1202
rect 802 1104 904 1208
rect -114 1026 904 1104
rect -114 1022 -12 1026
rect 802 1024 904 1026
<< via1 >>
rect 210 1768 302 1772
rect 210 1234 228 1768
rect 228 1234 280 1768
rect 280 1234 302 1768
rect 210 1230 302 1234
rect 494 1766 576 1772
rect 494 1234 508 1766
rect 508 1234 560 1766
rect 560 1234 576 1766
rect 494 1230 576 1234
<< metal2 >>
rect 200 1772 312 1802
rect 200 1230 210 1772
rect 302 1230 312 1772
rect 200 1202 312 1230
rect 480 1772 590 1800
rect 480 1230 494 1772
rect 576 1230 590 1772
rect 480 1202 590 1230
<< via2 >>
rect 210 1230 302 1772
rect 494 1230 576 1772
<< metal3 >>
rect 200 1772 312 1802
rect 200 1230 210 1772
rect 302 1230 312 1772
rect 200 818 312 1230
rect 480 1772 590 1800
rect 480 1230 494 1772
rect 576 1268 590 1772
rect 576 1230 592 1268
rect 480 832 592 1230
<< end >>
