magic
tech sky130A
magscale 1 2
timestamp 1698611618
<< error_p >>
rect -269 123 -211 129
rect -77 123 -19 129
rect 115 123 173 129
rect 307 123 365 129
rect -269 89 -257 123
rect -77 89 -65 123
rect 115 89 127 123
rect 307 89 319 123
rect -269 83 -211 89
rect -77 83 -19 89
rect 115 83 173 89
rect 307 83 365 89
rect -365 -89 -307 -83
rect -173 -89 -115 -83
rect 19 -89 77 -83
rect 211 -89 269 -83
rect -365 -123 -353 -89
rect -173 -123 -161 -89
rect 19 -123 31 -89
rect 211 -123 223 -89
rect -365 -129 -307 -123
rect -173 -129 -115 -123
rect 19 -129 77 -123
rect 211 -129 269 -123
<< nwell >>
rect -353 104 449 142
rect -449 -104 449 104
rect -449 -142 353 -104
<< pmos >>
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
<< pdiff >>
rect -413 30 -351 42
rect -413 -30 -401 30
rect -367 -30 -351 30
rect -413 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 413 42
rect 351 -30 367 30
rect 401 -30 413 30
rect 351 -42 413 -30
<< pdiffc >>
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
<< poly >>
rect -273 123 -207 139
rect -273 89 -257 123
rect -223 89 -207 123
rect -273 73 -207 89
rect -81 123 -15 139
rect -81 89 -65 123
rect -31 89 -15 123
rect -81 73 -15 89
rect 111 123 177 139
rect 111 89 127 123
rect 161 89 177 123
rect 111 73 177 89
rect 303 123 369 139
rect 303 89 319 123
rect 353 89 369 123
rect 303 73 369 89
rect -351 42 -321 68
rect -255 42 -225 73
rect -159 42 -129 68
rect -63 42 -33 73
rect 33 42 63 68
rect 129 42 159 73
rect 225 42 255 68
rect 321 42 351 73
rect -351 -73 -321 -42
rect -255 -68 -225 -42
rect -159 -73 -129 -42
rect -63 -68 -33 -42
rect 33 -73 63 -42
rect 129 -68 159 -42
rect 225 -73 255 -42
rect 321 -68 351 -42
rect -369 -89 -303 -73
rect -369 -123 -353 -89
rect -319 -123 -303 -89
rect -369 -139 -303 -123
rect -177 -89 -111 -73
rect -177 -123 -161 -89
rect -127 -123 -111 -89
rect -177 -139 -111 -123
rect 15 -89 81 -73
rect 15 -123 31 -89
rect 65 -123 81 -89
rect 15 -139 81 -123
rect 207 -89 273 -73
rect 207 -123 223 -89
rect 257 -123 273 -89
rect 207 -139 273 -123
<< polycont >>
rect -257 89 -223 123
rect -65 89 -31 123
rect 127 89 161 123
rect 319 89 353 123
rect -353 -123 -319 -89
rect -161 -123 -127 -89
rect 31 -123 65 -89
rect 223 -123 257 -89
<< locali >>
rect -273 89 -257 123
rect -223 89 -207 123
rect -81 89 -65 123
rect -31 89 -15 123
rect 111 89 127 123
rect 161 89 177 123
rect 303 89 319 123
rect 353 89 369 123
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect -369 -123 -353 -89
rect -319 -123 -303 -89
rect -177 -123 -161 -89
rect -127 -123 -111 -89
rect 15 -123 31 -89
rect 65 -123 81 -89
rect 207 -123 223 -89
rect 257 -123 273 -89
<< viali >>
rect -257 89 -223 123
rect -65 89 -31 123
rect 127 89 161 123
rect 319 89 353 123
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect -353 -123 -319 -89
rect -161 -123 -127 -89
rect 31 -123 65 -89
rect 223 -123 257 -89
<< metal1 >>
rect -269 123 -211 129
rect -269 89 -257 123
rect -223 89 -211 123
rect -269 83 -211 89
rect -77 123 -19 129
rect -77 89 -65 123
rect -31 89 -19 123
rect -77 83 -19 89
rect 115 123 173 129
rect 115 89 127 123
rect 161 89 173 123
rect 115 83 173 89
rect 307 123 365 129
rect 307 89 319 123
rect 353 89 365 123
rect 307 83 365 89
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect -365 -89 -307 -83
rect -365 -123 -353 -89
rect -319 -123 -307 -89
rect -365 -129 -307 -123
rect -173 -89 -115 -83
rect -173 -123 -161 -89
rect -127 -123 -115 -89
rect -173 -129 -115 -123
rect 19 -89 77 -83
rect 19 -123 31 -89
rect 65 -123 77 -89
rect 19 -129 77 -123
rect 211 -89 269 -83
rect 211 -123 223 -89
rect 257 -123 269 -89
rect 211 -129 269 -123
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
