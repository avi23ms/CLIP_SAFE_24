magic
tech sky130A
magscale 1 2
timestamp 1699103691
<< nwell >>
rect -929 104 1025 142
rect -1025 -104 1025 104
rect -1025 -142 929 -104
<< pmos >>
rect -927 -42 -897 42
rect -831 -42 -801 42
rect -735 -42 -705 42
rect -639 -42 -609 42
rect -543 -42 -513 42
rect -447 -42 -417 42
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
rect 417 -42 447 42
rect 513 -42 543 42
rect 609 -42 639 42
rect 705 -42 735 42
rect 801 -42 831 42
rect 897 -42 927 42
<< pdiff >>
rect -989 30 -927 42
rect -989 -30 -977 30
rect -943 -30 -927 30
rect -989 -42 -927 -30
rect -897 30 -831 42
rect -897 -30 -881 30
rect -847 -30 -831 30
rect -897 -42 -831 -30
rect -801 30 -735 42
rect -801 -30 -785 30
rect -751 -30 -735 30
rect -801 -42 -735 -30
rect -705 30 -639 42
rect -705 -30 -689 30
rect -655 -30 -639 30
rect -705 -42 -639 -30
rect -609 30 -543 42
rect -609 -30 -593 30
rect -559 -30 -543 30
rect -609 -42 -543 -30
rect -513 30 -447 42
rect -513 -30 -497 30
rect -463 -30 -447 30
rect -513 -42 -447 -30
rect -417 30 -351 42
rect -417 -30 -401 30
rect -367 -30 -351 30
rect -417 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 417 42
rect 351 -30 367 30
rect 401 -30 417 30
rect 351 -42 417 -30
rect 447 30 513 42
rect 447 -30 463 30
rect 497 -30 513 30
rect 447 -42 513 -30
rect 543 30 609 42
rect 543 -30 559 30
rect 593 -30 609 30
rect 543 -42 609 -30
rect 639 30 705 42
rect 639 -30 655 30
rect 689 -30 705 30
rect 639 -42 705 -30
rect 735 30 801 42
rect 735 -30 751 30
rect 785 -30 801 30
rect 735 -42 801 -30
rect 831 30 897 42
rect 831 -30 847 30
rect 881 -30 897 30
rect 831 -42 897 -30
rect 927 30 989 42
rect 927 -30 943 30
rect 977 -30 989 30
rect 927 -42 989 -30
<< pdiffc >>
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
<< poly >>
rect -849 123 -783 139
rect -849 89 -833 123
rect -799 89 -783 123
rect -849 73 -783 89
rect -657 123 -591 139
rect -657 89 -641 123
rect -607 89 -591 123
rect -657 73 -591 89
rect -465 123 -399 139
rect -465 89 -449 123
rect -415 89 -399 123
rect -465 73 -399 89
rect -273 123 -207 139
rect -273 89 -257 123
rect -223 89 -207 123
rect -273 73 -207 89
rect -81 123 -15 139
rect -81 89 -65 123
rect -31 89 -15 123
rect -81 73 -15 89
rect 111 123 177 139
rect 111 89 127 123
rect 161 89 177 123
rect 111 73 177 89
rect 303 123 369 139
rect 303 89 319 123
rect 353 89 369 123
rect 303 73 369 89
rect 495 123 561 139
rect 495 89 511 123
rect 545 89 561 123
rect 495 73 561 89
rect 687 123 753 139
rect 687 89 703 123
rect 737 89 753 123
rect 687 73 753 89
rect 879 123 945 139
rect 879 89 895 123
rect 929 89 945 123
rect 879 73 945 89
rect -927 42 -897 68
rect -831 42 -801 73
rect -735 42 -705 68
rect -639 42 -609 73
rect -543 42 -513 68
rect -447 42 -417 73
rect -351 42 -321 68
rect -255 42 -225 73
rect -159 42 -129 68
rect -63 42 -33 73
rect 33 42 63 68
rect 129 42 159 73
rect 225 42 255 68
rect 321 42 351 73
rect 417 42 447 68
rect 513 42 543 73
rect 609 42 639 68
rect 705 42 735 73
rect 801 42 831 68
rect 897 42 927 73
rect -927 -73 -897 -42
rect -831 -68 -801 -42
rect -735 -73 -705 -42
rect -639 -68 -609 -42
rect -543 -73 -513 -42
rect -447 -68 -417 -42
rect -351 -73 -321 -42
rect -255 -68 -225 -42
rect -159 -73 -129 -42
rect -63 -68 -33 -42
rect 33 -73 63 -42
rect 129 -68 159 -42
rect 225 -73 255 -42
rect 321 -68 351 -42
rect 417 -73 447 -42
rect 513 -68 543 -42
rect 609 -73 639 -42
rect 705 -68 735 -42
rect 801 -73 831 -42
rect 897 -68 927 -42
rect -945 -89 -879 -73
rect -945 -123 -929 -89
rect -895 -123 -879 -89
rect -945 -139 -879 -123
rect -753 -89 -687 -73
rect -753 -123 -737 -89
rect -703 -123 -687 -89
rect -753 -139 -687 -123
rect -561 -89 -495 -73
rect -561 -123 -545 -89
rect -511 -123 -495 -89
rect -561 -139 -495 -123
rect -369 -89 -303 -73
rect -369 -123 -353 -89
rect -319 -123 -303 -89
rect -369 -139 -303 -123
rect -177 -89 -111 -73
rect -177 -123 -161 -89
rect -127 -123 -111 -89
rect -177 -139 -111 -123
rect 15 -89 81 -73
rect 15 -123 31 -89
rect 65 -123 81 -89
rect 15 -139 81 -123
rect 207 -89 273 -73
rect 207 -123 223 -89
rect 257 -123 273 -89
rect 207 -139 273 -123
rect 399 -89 465 -73
rect 399 -123 415 -89
rect 449 -123 465 -89
rect 399 -139 465 -123
rect 591 -89 657 -73
rect 591 -123 607 -89
rect 641 -123 657 -89
rect 591 -139 657 -123
rect 783 -89 849 -73
rect 783 -123 799 -89
rect 833 -123 849 -89
rect 783 -139 849 -123
<< polycont >>
rect -833 89 -799 123
rect -641 89 -607 123
rect -449 89 -415 123
rect -257 89 -223 123
rect -65 89 -31 123
rect 127 89 161 123
rect 319 89 353 123
rect 511 89 545 123
rect 703 89 737 123
rect 895 89 929 123
rect -929 -123 -895 -89
rect -737 -123 -703 -89
rect -545 -123 -511 -89
rect -353 -123 -319 -89
rect -161 -123 -127 -89
rect 31 -123 65 -89
rect 223 -123 257 -89
rect 415 -123 449 -89
rect 607 -123 641 -89
rect 799 -123 833 -89
<< locali >>
rect -849 89 -833 123
rect -799 89 -783 123
rect -657 89 -641 123
rect -607 89 -591 123
rect -465 89 -449 123
rect -415 89 -399 123
rect -273 89 -257 123
rect -223 89 -207 123
rect -81 89 -65 123
rect -31 89 -15 123
rect 111 89 127 123
rect 161 89 177 123
rect 303 89 319 123
rect 353 89 369 123
rect 495 89 511 123
rect 545 89 561 123
rect 687 89 703 123
rect 737 89 753 123
rect 879 89 895 123
rect 929 89 945 123
rect -977 30 -943 46
rect -977 -46 -943 -30
rect -881 30 -847 46
rect -881 -46 -847 -30
rect -785 30 -751 46
rect -785 -46 -751 -30
rect -689 30 -655 46
rect -689 -46 -655 -30
rect -593 30 -559 46
rect -593 -46 -559 -30
rect -497 30 -463 46
rect -497 -46 -463 -30
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect 463 30 497 46
rect 463 -46 497 -30
rect 559 30 593 46
rect 559 -46 593 -30
rect 655 30 689 46
rect 655 -46 689 -30
rect 751 30 785 46
rect 751 -46 785 -30
rect 847 30 881 46
rect 847 -46 881 -30
rect 943 30 977 46
rect 943 -46 977 -30
rect -945 -123 -929 -89
rect -895 -123 -879 -89
rect -753 -123 -737 -89
rect -703 -123 -687 -89
rect -561 -123 -545 -89
rect -511 -123 -495 -89
rect -369 -123 -353 -89
rect -319 -123 -303 -89
rect -177 -123 -161 -89
rect -127 -123 -111 -89
rect 15 -123 31 -89
rect 65 -123 81 -89
rect 207 -123 223 -89
rect 257 -123 273 -89
rect 399 -123 415 -89
rect 449 -123 465 -89
rect 591 -123 607 -89
rect 641 -123 657 -89
rect 783 -123 799 -89
rect 833 -123 849 -89
<< viali >>
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
<< metal1 >>
rect -983 30 -937 42
rect -983 -30 -977 30
rect -943 -30 -937 30
rect -983 -42 -937 -30
rect -887 30 -841 42
rect -887 -30 -881 30
rect -847 -30 -841 30
rect -887 -42 -841 -30
rect -791 30 -745 42
rect -791 -30 -785 30
rect -751 -30 -745 30
rect -791 -42 -745 -30
rect -695 30 -649 42
rect -695 -30 -689 30
rect -655 -30 -649 30
rect -695 -42 -649 -30
rect -599 30 -553 42
rect -599 -30 -593 30
rect -559 -30 -553 30
rect -599 -42 -553 -30
rect -503 30 -457 42
rect -503 -30 -497 30
rect -463 -30 -457 30
rect -503 -42 -457 -30
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect 457 30 503 42
rect 457 -30 463 30
rect 497 -30 503 30
rect 457 -42 503 -30
rect 553 30 599 42
rect 553 -30 559 30
rect 593 -30 599 30
rect 553 -42 599 -30
rect 649 30 695 42
rect 649 -30 655 30
rect 689 -30 695 30
rect 649 -42 695 -30
rect 745 30 791 42
rect 745 -30 751 30
rect 785 -30 791 30
rect 745 -42 791 -30
rect 841 30 887 42
rect 841 -30 847 30
rect 881 -30 887 30
rect 841 -42 887 -30
rect 937 30 983 42
rect 937 -30 943 30
rect 977 -30 983 30
rect 937 -42 983 -30
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
