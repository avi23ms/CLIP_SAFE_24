magic
tech sky130A
magscale 1 2
timestamp 1698475453
<< error_s >>
rect 261 828 319 912
rect 349 828 407 912
rect 479 828 537 912
rect 567 828 625 912
rect 953 652 1015 736
rect 1045 652 1111 736
rect 1141 652 1207 736
rect 1237 652 1303 736
rect 1333 652 1399 736
rect 1429 652 1495 736
rect 1525 652 1591 736
rect 1621 652 1687 736
rect 1717 652 1783 736
rect 1813 652 1879 736
rect 1909 652 1975 736
rect 2005 652 2071 736
rect 2101 652 2167 736
rect 2197 652 2263 736
rect 2293 652 2359 736
rect 2389 652 2455 736
rect 2485 652 2551 736
rect 2581 652 2647 736
rect 2677 652 2743 736
rect 2773 652 2839 736
rect 2869 652 2935 736
rect 2965 652 3031 736
rect 3061 652 3127 736
rect 3157 652 3223 736
rect 3253 652 3319 736
rect 3349 652 3408 736
<< nwell >>
rect 228 1012 1238 1466
<< nsubdiff >>
rect 712 1340 854 1366
rect 712 1128 740 1340
rect 826 1128 854 1340
rect 712 1100 854 1128
<< nsubdiffcont >>
rect 740 1128 826 1340
<< locali >>
rect 712 1340 854 1366
rect 712 1128 740 1340
rect 826 1128 854 1340
rect 712 1100 854 1128
<< viali >>
rect 740 1128 826 1340
<< metal1 >>
rect 738 1368 862 1814
rect 712 1340 864 1368
rect 712 1128 740 1340
rect 826 1128 864 1340
rect 712 1100 864 1128
use capacitor_7  capacitor_7_0
timestamp 1698474969
transform 1 0 739 0 1 0
box -739 0 9807 2050
<< end >>
