magic
tech sky130A
magscale 1 2
timestamp 1698482903
<< metal1 >>
rect 12544 648 12578 824
rect 12416 -202 12864 -200
rect 12416 -256 12430 -202
rect 12836 -256 12864 -202
rect 12416 -262 12864 -256
rect 16560 -286 17248 -284
rect 12970 -288 23740 -286
rect 1334 -298 2508 -294
rect 4266 -298 5072 -292
rect 8048 -298 8662 -294
rect 1334 -300 10854 -298
rect 1334 -306 12234 -300
rect 1334 -492 1386 -306
rect 2462 -336 12234 -306
rect 2462 -338 10854 -336
rect 2464 -380 10854 -338
rect 2464 -472 4308 -380
rect 2462 -492 4308 -472
rect 1334 -516 4308 -492
rect 4266 -1608 4308 -516
rect 5016 -460 10854 -380
rect 5016 -516 8090 -460
rect 5016 -1608 5072 -516
rect 4266 -2310 5072 -1608
rect 8048 -1096 8090 -516
rect 8630 -516 10854 -460
rect 8630 -1096 8662 -516
rect 12198 -560 12234 -336
rect 12970 -302 23742 -288
rect 12970 -322 22496 -302
rect 12970 -560 13006 -322
rect 14427 -364 22496 -322
rect 14427 -508 21298 -364
rect 16560 -650 17248 -508
rect 16560 -844 16640 -650
rect 8048 -1852 8662 -1096
rect 16546 -1140 16640 -844
rect 17184 -844 17248 -650
rect 17184 -1140 17262 -844
rect 16546 -1196 17262 -1140
rect 21256 -1716 21298 -508
rect 21980 -490 22496 -364
rect 23662 -490 23742 -302
rect 21980 -502 23742 -490
rect 21980 -508 23176 -502
rect 21980 -1716 22030 -508
rect 21256 -2684 22030 -1716
<< via1 >>
rect 12430 -256 12836 -202
rect 1386 -338 2462 -306
rect 1386 -472 2464 -338
rect 1386 -492 2462 -472
rect 4308 -1608 5016 -380
rect 8090 -1096 8630 -460
rect 16640 -1140 17184 -650
rect 21298 -1716 21980 -364
rect 22496 -490 23662 -302
<< metal2 >>
rect 11778 15884 13440 15936
rect 11726 13798 13388 13850
rect 11892 11712 13380 11764
rect 11886 9626 13378 9678
rect 11938 7540 13314 7592
rect 11909 5456 13292 5508
rect 11886 3372 13244 3424
rect 11956 1284 13332 1336
rect 9818 -124 12354 -84
rect 1334 -306 2508 -294
rect 1334 -492 1386 -306
rect 2462 -338 2508 -306
rect 2464 -472 2508 -338
rect 2462 -492 2508 -472
rect 1334 -516 2508 -492
rect 4266 -380 5062 -298
rect 4266 -1608 4308 -380
rect 5016 -1608 5062 -380
rect 8044 -460 8670 -414
rect 8044 -1096 8090 -460
rect 8630 -1096 8670 -460
rect 8044 -1140 8670 -1096
rect 9818 -1110 9838 -124
rect 9916 -146 12354 -124
rect 9916 -1110 9942 -146
rect 12416 -202 12864 -200
rect 12416 -256 12430 -202
rect 12836 -222 12864 -202
rect 12836 -256 15842 -222
rect 12416 -262 15842 -256
rect 9818 -1138 9942 -1110
rect 15754 -290 15842 -262
rect 9835 -1585 9897 -1138
rect 15754 -1140 15774 -290
rect 15830 -1140 15842 -290
rect 21236 -364 22030 -282
rect 16560 -650 17258 -566
rect 16560 -844 16640 -650
rect 15754 -1174 15842 -1140
rect 16546 -1140 16640 -844
rect 17184 -844 17258 -650
rect 17184 -1140 17262 -844
rect 16546 -1196 17262 -1140
rect 4266 -1690 5062 -1608
rect 21236 -1716 21298 -364
rect 21980 -1716 22030 -364
rect 22452 -302 23742 -288
rect 22452 -490 22496 -302
rect 23662 -490 23742 -302
rect 22452 -502 23742 -490
rect 21236 -1860 22030 -1716
<< via2 >>
rect 1386 -338 2462 -306
rect 1386 -472 2464 -338
rect 1386 -492 2462 -472
rect 4308 -1608 5016 -380
rect 8090 -1096 8630 -460
rect 9838 -1110 9916 -124
rect 15774 -1140 15830 -290
rect 16640 -1140 17184 -650
rect 21298 -1716 21980 -364
rect 22496 -490 23662 -302
<< metal3 >>
rect 12910 15813 13417 15815
rect 11658 15805 12314 15806
rect 11658 15542 12400 15805
rect 11874 13734 12400 15542
rect 11674 13488 12400 13734
rect 11874 11648 12400 13488
rect 11699 11402 12400 11648
rect 11874 9562 12400 11402
rect 11689 9316 12400 9562
rect 11874 7476 12400 9316
rect 11755 7230 12400 7476
rect 11874 5392 12400 7230
rect 11724 5146 12400 5392
rect 11874 3308 12400 5146
rect 11741 3062 12400 3308
rect 11874 1224 12400 3062
rect 11782 960 12400 1224
rect 12718 15573 13417 15813
rect 12718 13724 13244 15573
rect 12718 13478 13477 13724
rect 12718 11638 13244 13478
rect 12718 11392 13403 11638
rect 12718 9552 13244 11392
rect 12718 9306 13389 9552
rect 12718 7466 13244 9306
rect 12718 7220 13407 7466
rect 12718 5382 13244 7220
rect 12718 5136 13455 5382
rect 1338 -294 1428 167
rect 12272 112 12336 960
rect 12718 942 13244 5136
rect 5916 -10 12336 112
rect 1334 -306 2508 -294
rect 1334 -492 1386 -306
rect 2462 -338 2508 -306
rect 2464 -472 2508 -338
rect 2462 -492 2508 -472
rect 1334 -516 2508 -492
rect 4266 -380 5062 -298
rect 1338 -519 1428 -516
rect 4266 -1608 4308 -380
rect 5016 -1608 5062 -380
rect 4266 -1690 5062 -1608
rect 5916 -2614 6130 -10
rect 12272 -74 12336 -10
rect 12792 98 12856 942
rect 12792 95 20200 98
rect 12792 -36 20312 95
rect 9818 -124 9942 -84
rect 12799 -95 20312 -36
rect 8044 -460 8670 -414
rect 8044 -1096 8090 -460
rect 8630 -1096 8670 -460
rect 8044 -1140 8670 -1096
rect 9818 -1110 9838 -124
rect 9916 -1110 9942 -124
rect 15754 -290 15842 -222
rect 15754 -550 15774 -290
rect 9818 -1138 9942 -1110
rect 15748 -1140 15774 -550
rect 15830 -550 15842 -290
rect 15830 -1140 15846 -550
rect 16558 -552 17258 -520
rect 16558 -650 17268 -552
rect 16558 -844 16640 -650
rect 16546 -1140 16640 -844
rect 17184 -1140 17268 -650
rect 15754 -1174 15842 -1140
rect 15756 -1474 15832 -1174
rect 16546 -1196 17262 -1140
rect 16558 -1226 17258 -1196
rect 20122 -2396 20312 -95
rect 21236 -364 22030 -282
rect 23655 -288 23745 119
rect 21236 -1716 21298 -364
rect 21980 -1716 22030 -364
rect 22452 -302 23745 -288
rect 22452 -490 22496 -302
rect 23662 -490 23745 -302
rect 22452 -502 23745 -490
rect 23655 -503 23745 -502
rect 21236 -1860 22030 -1716
rect 12446 -6994 12518 -6620
<< via3 >>
rect 4308 -1608 5016 -380
rect 8090 -1096 8630 -460
rect 16640 -1140 17184 -650
rect 21298 -1716 21980 -364
<< metal4 >>
rect 667 -5056 1235 568
rect 4266 -380 5072 -292
rect 4266 -1608 4308 -380
rect 5016 -1608 5072 -380
rect 4266 -2310 5072 -1608
rect 8048 -460 8662 -294
rect 8048 -1096 8090 -460
rect 8630 -1096 8662 -460
rect 21256 -364 22030 -286
rect 8048 -1852 8662 -1096
rect 16574 -650 17254 -574
rect 16574 -1140 16640 -650
rect 17184 -1140 17254 -650
rect 16574 -1408 17254 -1140
rect 21256 -1716 21298 -364
rect 21980 -1716 22030 -364
rect 21256 -2684 22030 -1716
rect 667 -5624 11584 -5056
<< metal5 >>
rect 24493 -4695 25083 585
rect 13677 -5285 25083 -4695
use capacitors_8  capacitors_8_0 ~/Desktop/charge_pumps2/layout_files2
timestamp 1698479562
transform 1 0 1291 0 1 14846
box -1291 -14846 10740 2058
use capacitors_8  capacitors_8_1
timestamp 1698479562
transform -1 0 23792 0 1 14836
box -1291 -14846 10740 2058
use clock  clock_0 ~/Desktop/charge_pumps2/layout_files2
timestamp 1698410772
transform 0 -1 12414 1 0 -6496
box -410 -1832 6030 1274
use pmos_cp1  pmos_cp1_0 ~/Desktop/charge_pumps2/layout_files2
timestamp 1698464655
transform 1 0 12252 0 1 -82
box -14 -278 858 754
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_0
timestamp 0
transform -1 0 16844 0 1 -2266
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_1
timestamp 0
transform 1 0 8830 0 1 -2176
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_2
timestamp 0
transform 1 0 5052 0 1 -2796
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_3
timestamp 0
transform -1 0 21206 0 1 -3076
box -1086 -940 1086 940
<< labels >>
rlabel metal1 12552 772 12552 772 1 out
port 30 n
rlabel metal1 11752 -322 11752 -322 1 clk
port 31 n
rlabel metal1 13296 -304 13296 -302 1 clkb
port 32 n
rlabel metal3 12474 -6950 12474 -6950 1 clk_in
port 33 n
rlabel metal3 12088 15446 12088 15446 1 input1
port 34 n
rlabel metal3 12964 15418 12964 15418 1 input2
port 35 n
rlabel space 166 8424 166 8424 1 vdd
port 36 n
rlabel space 810 9748 810 9748 1 gnd
port 37 n
rlabel metal4 862 -3106 862 -3106 1 vdd
port 38 n
rlabel metal5 18556 -5038 18556 -5038 1 gnd
port 39 n
<< end >>
