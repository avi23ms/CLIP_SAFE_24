magic
tech sky130A
magscale 1 2
timestamp 1697921677
<< metal1 >>
rect 150 1513 312 1583
rect 3226 1550 3236 1614
rect 3334 1550 3344 1614
rect 1878 982 1976 986
rect 1878 914 1914 982
rect 1986 914 1996 982
rect 1878 902 1976 914
rect 477 656 582 659
rect 470 604 480 656
rect 564 604 582 656
rect 477 577 582 604
rect 270 78 312 442
rect 412 336 486 360
rect 412 320 494 336
rect 412 282 500 320
rect 420 258 500 282
rect 464 256 500 258
rect 464 214 1600 256
rect 464 206 500 214
rect 770 -129 813 -59
rect 2714 -66 2724 -42
rect 2498 -114 2724 -66
rect 2714 -124 2724 -114
rect 2788 -124 2798 -42
rect 1794 -1028 1804 -966
rect 1886 -1028 1896 -966
rect 2852 -1077 2901 494
rect 2491 -1126 2901 -1077
<< via1 >>
rect 3236 1550 3334 1614
rect 1914 914 1986 982
rect 480 604 564 656
rect 2724 -124 2788 -42
rect 1804 -1028 1886 -966
<< metal2 >>
rect 3236 1614 3334 1624
rect 3334 1556 3660 1611
rect 3236 1540 3334 1550
rect 1914 982 1986 992
rect 1986 924 2636 972
rect 1914 904 1986 914
rect 480 656 564 666
rect 480 594 564 604
rect 492 -1008 532 594
rect 880 14 920 872
rect 880 -26 1724 14
rect 1684 -924 1724 -26
rect 464 -1117 532 -1008
rect 1804 -966 1886 -956
rect 2588 -974 2636 924
rect 2724 -42 2788 -32
rect 3605 -54 3660 1556
rect 2788 -106 3660 -54
rect 3605 -107 3660 -106
rect 2724 -134 2788 -124
rect 1886 -1014 2636 -974
rect 2588 -1018 2636 -1014
rect 1804 -1038 1886 -1028
rect 464 -1120 510 -1117
use cmfb  cmfb_0
timestamp 1697921677
transform 1 0 -54 0 1 -439
box 203 439 3639 2056
use integrator2  integrator2_0
timestamp 1697921677
transform 1 0 -1633 0 1 -3755
box 1247 441 5619 3693
use sky130_fd_pr__nfet_01v8_TABC9M  sky130_fd_pr__nfet_01v8_TABC9M_0
timestamp 1697388782
transform -1 0 396 0 -1 176
box -246 -310 246 310
<< labels >>
rlabel metal1 2761 -1077 2761 -1077 1 gnd
rlabel metal2 916 91 916 91 3 vo2
rlabel metal1 1072 256 1072 256 1 Vbias
rlabel metal2 2538 -977 2538 -976 1 Vbn
<< end >>
