magic
tech sky130A
magscale 1 2
timestamp 1698651669
<< error_s >>
rect 4606 1913 5584 1942
rect 4568 1875 5546 1904
rect 4824 1842 4964 1869
rect 4846 1831 4882 1832
rect 4846 1804 4926 1831
rect 4846 1794 4882 1804
rect 4744 1777 4792 1794
rect 4822 1778 4882 1794
rect 4812 1777 4882 1778
rect 4744 1749 4792 1766
rect 4812 1743 4828 1777
rect 4846 1761 4882 1777
rect 4732 1724 4828 1743
rect 4708 1717 4828 1724
rect 4674 1706 4828 1717
rect 4708 1693 4828 1706
rect 4732 1690 4828 1693
rect 4702 1678 4710 1689
rect 4732 1677 4754 1689
rect 4710 1672 4754 1677
rect 4732 1665 4754 1672
rect 4696 1644 4711 1659
rect 4696 1618 4754 1644
rect 4708 1501 4742 1618
rect 5441 1606 5486 1617
rect 5452 1489 5486 1606
rect 5496 1524 5540 1547
rect 5496 1489 5498 1524
rect 5440 1442 5498 1489
rect 4770 1418 5498 1442
rect 5524 1496 5540 1519
rect 5524 1476 5526 1496
rect 4770 1408 5462 1409
rect 4758 1402 5410 1405
rect 5524 1389 5652 1476
rect 4730 1374 5410 1377
rect 4732 1370 5424 1371
rect 4546 1318 5538 1355
rect 4682 990 4697 1005
rect 4682 964 4740 990
rect 4694 847 4728 964
rect 5427 952 5472 963
rect 5438 835 5472 952
rect 5778 941 5892 1222
rect 5930 1180 5945 1195
rect 5960 1192 5982 1225
rect 5952 1180 5982 1192
rect 5930 1154 5982 1180
rect 5988 1158 6010 1253
rect 5942 1037 5976 1154
rect 5952 1021 5976 1037
rect 5986 1153 6010 1158
rect 5986 1025 6020 1153
rect 6058 1038 6146 1064
rect 6226 1038 6262 1064
rect 6058 1035 6262 1038
rect 6058 1025 6146 1035
rect 5986 1013 6032 1025
rect 6100 1021 6134 1025
rect 5957 992 6032 1013
rect 5957 978 6038 992
rect 6112 989 6168 1010
rect 6172 1007 6208 1010
rect 6084 987 6168 989
rect 6084 978 6122 987
rect 5957 966 6032 978
rect 5974 954 6032 966
rect 6078 964 6122 978
rect 6078 961 6088 964
rect 6112 961 6122 964
rect 5988 941 6016 954
rect 6078 944 6122 961
rect 6192 959 6208 1007
rect 6226 993 6262 1035
rect 5778 934 6016 941
rect 6084 936 6122 944
rect 5544 931 5546 934
rect 5592 931 6016 934
rect 5778 913 5892 931
rect 5984 929 6016 931
rect 5988 928 6016 929
rect 6112 922 6122 936
rect 5778 906 5970 913
rect 5516 903 5546 906
rect 5592 903 5970 906
rect 5778 846 5892 903
rect 5958 901 5970 903
rect 5426 788 5484 835
rect 4756 764 5484 788
rect 4756 754 5448 755
rect 4752 748 5450 751
rect 4752 743 4768 748
rect 4752 720 5422 723
rect 4752 717 4796 720
rect 4718 716 5410 717
rect 4752 715 4796 716
rect 4652 672 4654 677
rect 4680 644 4682 677
rect 5472 587 5488 638
rect 5506 621 5542 692
rect 4622 553 5644 569
rect 4618 498 5644 553
rect 4508 482 5644 498
rect 4504 410 5644 482
rect 4508 301 5644 410
rect 4508 230 5530 301
use comparator_final_compact  comparator_final_compact_0
timestamp 1698651669
transform 1 0 6806 0 1 2474
box -2212 -2214 6449 1614
use integrator_full_new_compact  integrator_full_new_compact_0
timestamp 1698651669
transform 1 0 386 0 1 3329
box -386 -3329 4003 1133
use reference  reference_0
timestamp 1698586885
transform 1 0 4546 0 1 1318
box -66 -1120 1956 620
<< end >>
