magic
tech sky130A
timestamp 1726930802
<< error_p >>
rect 31 41 48 44
rect 31 -41 34 41
rect 45 -41 48 41
rect 31 -44 48 -41
<< nmos >>
rect -25 -50 25 50
<< ndiff >>
rect -54 44 -25 50
rect -54 -44 -48 44
rect -31 -44 -25 44
rect -54 -50 -25 -44
rect 25 -50 54 50
<< ndiffc >>
rect -48 -44 -31 44
<< poly >>
rect -25 50 25 63
rect -25 -63 25 -50
<< locali >>
rect -48 44 -31 52
rect -48 -52 -31 -44
<< viali >>
rect -48 -44 -31 44
rect 31 -44 48 44
<< metal1 >>
rect -51 44 -28 50
rect -51 -44 -48 44
rect -31 -44 -28 44
rect -51 -50 -28 -44
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
