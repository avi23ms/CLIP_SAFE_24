magic
tech sky130A
magscale 1 2
timestamp 1727421560
<< viali >>
rect 5365 10217 5399 10251
rect 5917 10217 5951 10251
rect 1409 10013 1443 10047
rect 5181 10013 5215 10047
rect 5641 9945 5675 9979
rect 1593 9877 1627 9911
rect 5365 9673 5399 9707
rect 5549 9605 5583 9639
rect 5733 9605 5767 9639
rect 1501 9537 1535 9571
rect 3801 9537 3835 9571
rect 5181 9537 5215 9571
rect 5457 9537 5491 9571
rect 5917 9537 5951 9571
rect 3709 9469 3743 9503
rect 5733 9401 5767 9435
rect 1777 9333 1811 9367
rect 3433 9333 3467 9367
rect 3801 9333 3835 9367
rect 6101 9333 6135 9367
rect 5825 9061 5859 9095
rect 3341 8993 3375 9027
rect 4169 8993 4203 9027
rect 5457 8993 5491 9027
rect 5549 8993 5583 9027
rect 3433 8925 3467 8959
rect 3525 8925 3559 8959
rect 4077 8925 4111 8959
rect 4261 8925 4295 8959
rect 5733 8925 5767 8959
rect 5917 8925 5951 8959
rect 6009 8925 6043 8959
rect 6193 8925 6227 8959
rect 3157 8789 3191 8823
rect 3893 8789 3927 8823
rect 4813 8789 4847 8823
rect 6193 8585 6227 8619
rect 4353 8449 4387 8483
rect 4445 8381 4479 8415
rect 4721 8381 4755 8415
rect 3065 8245 3099 8279
rect 5917 8041 5951 8075
rect 3341 7905 3375 7939
rect 4169 7905 4203 7939
rect 3065 7769 3099 7803
rect 4445 7769 4479 7803
rect 1593 7701 1627 7735
rect 4537 7497 4571 7531
rect 6193 7497 6227 7531
rect 3157 7361 3191 7395
rect 3433 7361 3467 7395
rect 3709 7361 3743 7395
rect 4077 7361 4111 7395
rect 4353 7361 4387 7395
rect 4813 7361 4847 7395
rect 5641 7361 5675 7395
rect 2881 7293 2915 7327
rect 3249 7293 3283 7327
rect 5089 7293 5123 7327
rect 3525 7225 3559 7259
rect 3617 7225 3651 7259
rect 4169 7225 4203 7259
rect 4261 7225 4295 7259
rect 4629 7225 4663 7259
rect 1409 7157 1443 7191
rect 4997 7157 5031 7191
rect 2605 6953 2639 6987
rect 3249 6953 3283 6987
rect 3801 6953 3835 6987
rect 4353 6953 4387 6987
rect 4537 6953 4571 6987
rect 2513 6817 2547 6851
rect 2881 6817 2915 6851
rect 2973 6817 3007 6851
rect 4077 6817 4111 6851
rect 4169 6817 4203 6851
rect 6101 6817 6135 6851
rect 1593 6749 1627 6783
rect 1869 6749 1903 6783
rect 2053 6749 2087 6783
rect 2145 6749 2179 6783
rect 2329 6749 2363 6783
rect 2789 6749 2823 6783
rect 3065 6749 3099 6783
rect 3249 6749 3283 6783
rect 3341 6749 3375 6783
rect 3985 6749 4019 6783
rect 4629 6749 4663 6783
rect 4721 6749 4755 6783
rect 5825 6749 5859 6783
rect 1961 6681 1995 6715
rect 3617 6613 3651 6647
rect 1593 6409 1627 6443
rect 5089 6409 5123 6443
rect 1409 6273 1443 6307
rect 2605 6273 2639 6307
rect 3065 6273 3099 6307
rect 4905 6273 4939 6307
rect 5917 6273 5951 6307
rect 2789 6137 2823 6171
rect 4353 6069 4387 6103
rect 6101 6069 6135 6103
rect 3801 5865 3835 5899
rect 4169 5865 4203 5899
rect 4905 5729 4939 5763
rect 4997 5729 5031 5763
rect 5107 5729 5141 5763
rect 1409 5661 1443 5695
rect 3985 5661 4019 5695
rect 4261 5661 4295 5695
rect 5825 5593 5859 5627
rect 1593 5525 1627 5559
rect 4721 5525 4755 5559
rect 6101 5525 6135 5559
rect 2053 5253 2087 5287
rect 3249 5185 3283 5219
rect 3525 5185 3559 5219
rect 4169 5185 4203 5219
rect 4641 5185 4675 5219
rect 4813 5185 4847 5219
rect 4905 5185 4939 5219
rect 5273 5185 5307 5219
rect 6009 5185 6043 5219
rect 2513 5117 2547 5151
rect 2605 5117 2639 5151
rect 2973 5117 3007 5151
rect 3893 5117 3927 5151
rect 3985 5117 4019 5151
rect 4721 5117 4755 5151
rect 5089 5117 5123 5151
rect 5549 5117 5583 5151
rect 5917 5117 5951 5151
rect 2053 5049 2087 5083
rect 3065 5049 3099 5083
rect 3709 5049 3743 5083
rect 4353 5049 4387 5083
rect 5641 5049 5675 5083
rect 2789 4981 2823 5015
rect 3433 4981 3467 5015
rect 4445 4981 4479 5015
rect 5457 4981 5491 5015
rect 6009 4981 6043 5015
rect 3893 4641 3927 4675
rect 4077 4641 4111 4675
rect 4629 4641 4663 4675
rect 2099 4573 2133 4607
rect 2484 4573 2518 4607
rect 2605 4573 2639 4607
rect 3249 4573 3283 4607
rect 3985 4573 4019 4607
rect 4353 4573 4387 4607
rect 2237 4505 2271 4539
rect 2329 4505 2363 4539
rect 2697 4505 2731 4539
rect 1961 4437 1995 4471
rect 4261 4437 4295 4471
rect 6101 4437 6135 4471
rect 3525 4097 3559 4131
rect 3801 4097 3835 4131
rect 1501 4029 1535 4063
rect 1777 4029 1811 4063
rect 3617 4029 3651 4063
rect 4353 4029 4387 4063
rect 4629 4029 4663 4063
rect 3249 3961 3283 3995
rect 3709 3961 3743 3995
rect 3341 3893 3375 3927
rect 6101 3893 6135 3927
rect 5089 3689 5123 3723
rect 5641 3689 5675 3723
rect 5825 3689 5859 3723
rect 3341 3553 3375 3587
rect 5917 3553 5951 3587
rect 3801 3485 3835 3519
rect 6009 3485 6043 3519
rect 3065 3417 3099 3451
rect 1593 3349 1627 3383
rect 3433 3145 3467 3179
rect 3801 3145 3835 3179
rect 4353 3145 4387 3179
rect 6101 3145 6135 3179
rect 1409 3009 1443 3043
rect 3065 3009 3099 3043
rect 3249 3009 3283 3043
rect 3985 3009 4019 3043
rect 4077 3009 4111 3043
rect 4169 3009 4203 3043
rect 4537 3009 4571 3043
rect 4849 3009 4883 3043
rect 5917 3009 5951 3043
rect 1685 2941 1719 2975
rect 4721 2941 4755 2975
rect 4629 2873 4663 2907
rect 3065 2805 3099 2839
rect 5365 2397 5399 2431
rect 5825 2329 5859 2363
rect 5549 2261 5583 2295
rect 6101 2261 6135 2295
<< metal1 >>
rect 1104 10362 6532 10384
rect 1104 10310 1628 10362
rect 1680 10310 1692 10362
rect 1744 10310 1756 10362
rect 1808 10310 1820 10362
rect 1872 10310 1884 10362
rect 1936 10310 2984 10362
rect 3036 10310 3048 10362
rect 3100 10310 3112 10362
rect 3164 10310 3176 10362
rect 3228 10310 3240 10362
rect 3292 10310 4340 10362
rect 4392 10310 4404 10362
rect 4456 10310 4468 10362
rect 4520 10310 4532 10362
rect 4584 10310 4596 10362
rect 4648 10310 5696 10362
rect 5748 10310 5760 10362
rect 5812 10310 5824 10362
rect 5876 10310 5888 10362
rect 5940 10310 5952 10362
rect 6004 10310 6532 10362
rect 1104 10288 6532 10310
rect 5350 10208 5356 10260
rect 5408 10208 5414 10260
rect 5905 10251 5963 10257
rect 5905 10217 5917 10251
rect 5951 10248 5963 10251
rect 6362 10248 6368 10260
rect 5951 10220 6368 10248
rect 5951 10217 5963 10220
rect 5905 10211 5963 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 934 10004 940 10056
rect 992 10044 998 10056
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 992 10016 1409 10044
rect 992 10004 998 10016
rect 1397 10013 1409 10016
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 5442 10044 5448 10056
rect 5215 10016 5448 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 5629 9979 5687 9985
rect 5629 9976 5641 9979
rect 5408 9948 5641 9976
rect 5408 9936 5414 9948
rect 5629 9945 5641 9948
rect 5675 9945 5687 9979
rect 5629 9939 5687 9945
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 3510 9908 3516 9920
rect 1627 9880 3516 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 3510 9868 3516 9880
rect 3568 9868 3574 9920
rect 1104 9818 6670 9840
rect 1104 9766 2288 9818
rect 2340 9766 2352 9818
rect 2404 9766 2416 9818
rect 2468 9766 2480 9818
rect 2532 9766 2544 9818
rect 2596 9766 3644 9818
rect 3696 9766 3708 9818
rect 3760 9766 3772 9818
rect 3824 9766 3836 9818
rect 3888 9766 3900 9818
rect 3952 9766 5000 9818
rect 5052 9766 5064 9818
rect 5116 9766 5128 9818
rect 5180 9766 5192 9818
rect 5244 9766 5256 9818
rect 5308 9766 6356 9818
rect 6408 9766 6420 9818
rect 6472 9766 6484 9818
rect 6536 9766 6548 9818
rect 6600 9766 6612 9818
rect 6664 9766 6670 9818
rect 1104 9744 6670 9766
rect 5350 9664 5356 9716
rect 5408 9664 5414 9716
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 5537 9639 5595 9645
rect 4304 9608 5488 9636
rect 4304 9596 4310 9608
rect 934 9528 940 9580
rect 992 9568 998 9580
rect 1489 9571 1547 9577
rect 1489 9568 1501 9571
rect 992 9540 1501 9568
rect 992 9528 998 9540
rect 1489 9537 1501 9540
rect 1535 9537 1547 9571
rect 1489 9531 1547 9537
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 5460 9577 5488 9608
rect 5537 9605 5549 9639
rect 5583 9636 5595 9639
rect 5721 9639 5779 9645
rect 5583 9608 5672 9636
rect 5583 9605 5595 9608
rect 5537 9599 5595 9605
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 2740 9540 3801 9568
rect 2740 9528 2746 9540
rect 3789 9537 3801 9540
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5445 9571 5503 9577
rect 5215 9540 5396 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5368 9512 5396 9540
rect 5445 9537 5457 9571
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 3697 9503 3755 9509
rect 3697 9469 3709 9503
rect 3743 9500 3755 9503
rect 4890 9500 4896 9512
rect 3743 9472 4896 9500
rect 3743 9469 3755 9472
rect 3697 9463 3755 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5350 9460 5356 9512
rect 5408 9460 5414 9512
rect 5644 9432 5672 9608
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 6086 9636 6092 9648
rect 5767 9608 6092 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 6086 9596 6092 9608
rect 6144 9596 6150 9648
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 6270 9568 6276 9580
rect 5951 9540 6276 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 5460 9404 5672 9432
rect 5721 9435 5779 9441
rect 5460 9376 5488 9404
rect 5721 9401 5733 9435
rect 5767 9432 5779 9435
rect 6178 9432 6184 9444
rect 5767 9404 6184 9432
rect 5767 9401 5779 9404
rect 5721 9395 5779 9401
rect 6178 9392 6184 9404
rect 6236 9392 6242 9444
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 1946 9364 1952 9376
rect 1811 9336 1952 9364
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 3418 9324 3424 9376
rect 3476 9324 3482 9376
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3568 9336 3801 9364
rect 3568 9324 3574 9336
rect 3789 9333 3801 9336
rect 3835 9364 3847 9367
rect 5442 9364 5448 9376
rect 3835 9336 5448 9364
rect 3835 9333 3847 9336
rect 3789 9327 3847 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 6089 9367 6147 9373
rect 6089 9333 6101 9367
rect 6135 9364 6147 9367
rect 6730 9364 6736 9376
rect 6135 9336 6736 9364
rect 6135 9333 6147 9336
rect 6089 9327 6147 9333
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 1104 9274 6532 9296
rect 1104 9222 1628 9274
rect 1680 9222 1692 9274
rect 1744 9222 1756 9274
rect 1808 9222 1820 9274
rect 1872 9222 1884 9274
rect 1936 9222 2984 9274
rect 3036 9222 3048 9274
rect 3100 9222 3112 9274
rect 3164 9222 3176 9274
rect 3228 9222 3240 9274
rect 3292 9222 4340 9274
rect 4392 9222 4404 9274
rect 4456 9222 4468 9274
rect 4520 9222 4532 9274
rect 4584 9222 4596 9274
rect 4648 9222 5696 9274
rect 5748 9222 5760 9274
rect 5812 9222 5824 9274
rect 5876 9222 5888 9274
rect 5940 9222 5952 9274
rect 6004 9222 6532 9274
rect 1104 9200 6532 9222
rect 5442 9120 5448 9172
rect 5500 9120 5506 9172
rect 4246 9092 4252 9104
rect 4080 9064 4252 9092
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 9024 3387 9027
rect 4080 9024 4108 9064
rect 4246 9052 4252 9064
rect 4304 9052 4310 9104
rect 5460 9092 5488 9120
rect 5813 9095 5871 9101
rect 5813 9092 5825 9095
rect 5460 9064 5825 9092
rect 5813 9061 5825 9064
rect 5859 9061 5871 9095
rect 5813 9055 5871 9061
rect 6086 9052 6092 9104
rect 6144 9052 6150 9104
rect 6178 9052 6184 9104
rect 6236 9052 6242 9104
rect 3375 8996 4108 9024
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 4080 8968 4108 8996
rect 4157 9027 4215 9033
rect 4157 8993 4169 9027
rect 4203 9024 4215 9027
rect 4706 9024 4712 9036
rect 4203 8996 4712 9024
rect 4203 8993 4215 8996
rect 4157 8987 4215 8993
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 3436 8888 3464 8919
rect 3510 8916 3516 8968
rect 3568 8916 3574 8968
rect 4062 8916 4068 8968
rect 4120 8916 4126 8968
rect 4172 8888 4200 8987
rect 4706 8984 4712 8996
rect 4764 9024 4770 9036
rect 5445 9027 5503 9033
rect 4764 8996 5396 9024
rect 4764 8984 4770 8996
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8958 4307 8959
rect 4295 8956 4384 8958
rect 5368 8956 5396 8996
rect 5445 8993 5457 9027
rect 5491 9024 5503 9027
rect 5537 9027 5595 9033
rect 5537 9024 5549 9027
rect 5491 8996 5549 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 5537 8993 5549 8996
rect 5583 8993 5595 9027
rect 6104 9024 6132 9052
rect 5537 8987 5595 8993
rect 5736 8996 6132 9024
rect 5736 8965 5764 8996
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 4295 8930 5304 8956
rect 4295 8925 4307 8930
rect 4356 8928 5304 8930
rect 5368 8928 5733 8956
rect 4249 8919 4307 8925
rect 3436 8860 4200 8888
rect 5276 8888 5304 8928
rect 5721 8925 5733 8928
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6086 8956 6092 8968
rect 6043 8928 6092 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 5350 8888 5356 8900
rect 5276 8860 5356 8888
rect 5350 8848 5356 8860
rect 5408 8888 5414 8900
rect 5920 8888 5948 8919
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6196 8965 6224 9052
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8925 6239 8959
rect 6181 8919 6239 8925
rect 5408 8860 6776 8888
rect 5408 8848 5414 8860
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 3145 8823 3203 8829
rect 3145 8820 3157 8823
rect 2924 8792 3157 8820
rect 2924 8780 2930 8792
rect 3145 8789 3157 8792
rect 3191 8789 3203 8823
rect 3145 8783 3203 8789
rect 3881 8823 3939 8829
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 4246 8820 4252 8832
rect 3927 8792 4252 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4798 8780 4804 8832
rect 4856 8780 4862 8832
rect 1104 8730 6670 8752
rect 1104 8678 2288 8730
rect 2340 8678 2352 8730
rect 2404 8678 2416 8730
rect 2468 8678 2480 8730
rect 2532 8678 2544 8730
rect 2596 8678 3644 8730
rect 3696 8678 3708 8730
rect 3760 8678 3772 8730
rect 3824 8678 3836 8730
rect 3888 8678 3900 8730
rect 3952 8678 5000 8730
rect 5052 8678 5064 8730
rect 5116 8678 5128 8730
rect 5180 8678 5192 8730
rect 5244 8678 5256 8730
rect 5308 8678 6356 8730
rect 6408 8678 6420 8730
rect 6472 8678 6484 8730
rect 6536 8678 6548 8730
rect 6600 8678 6612 8730
rect 6664 8678 6670 8730
rect 1104 8656 6670 8678
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 6748 8616 6776 8860
rect 6227 8588 6776 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 1946 8508 1952 8560
rect 2004 8548 2010 8560
rect 4982 8548 4988 8560
rect 2004 8520 4988 8548
rect 2004 8508 2010 8520
rect 4982 8508 4988 8520
rect 5040 8548 5046 8560
rect 5040 8520 5198 8548
rect 5040 8508 5046 8520
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 4212 8452 4353 8480
rect 4212 8440 4218 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4433 8415 4491 8421
rect 4433 8412 4445 8415
rect 3344 8384 4445 8412
rect 3344 8288 3372 8384
rect 4433 8381 4445 8384
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 4798 8412 4804 8424
rect 4755 8384 4804 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 3053 8279 3111 8285
rect 3053 8245 3065 8279
rect 3099 8276 3111 8279
rect 3326 8276 3332 8288
rect 3099 8248 3332 8276
rect 3099 8245 3111 8248
rect 3053 8239 3111 8245
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 1104 8186 6532 8208
rect 1104 8134 1628 8186
rect 1680 8134 1692 8186
rect 1744 8134 1756 8186
rect 1808 8134 1820 8186
rect 1872 8134 1884 8186
rect 1936 8134 2984 8186
rect 3036 8134 3048 8186
rect 3100 8134 3112 8186
rect 3164 8134 3176 8186
rect 3228 8134 3240 8186
rect 3292 8134 4340 8186
rect 4392 8134 4404 8186
rect 4456 8134 4468 8186
rect 4520 8134 4532 8186
rect 4584 8134 4596 8186
rect 4648 8134 5696 8186
rect 5748 8134 5760 8186
rect 5812 8134 5824 8186
rect 5876 8134 5888 8186
rect 5940 8134 5952 8186
rect 6004 8134 6532 8186
rect 1104 8112 6532 8134
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 3510 8072 3516 8084
rect 3292 8044 3516 8072
rect 3292 8032 3298 8044
rect 3510 8032 3516 8044
rect 3568 8072 3574 8084
rect 5626 8072 5632 8084
rect 3568 8044 5632 8072
rect 3568 8032 3574 8044
rect 5626 8032 5632 8044
rect 5684 8072 5690 8084
rect 5905 8075 5963 8081
rect 5905 8072 5917 8075
rect 5684 8044 5917 8072
rect 5684 8032 5690 8044
rect 5905 8041 5917 8044
rect 5951 8072 5963 8075
rect 6270 8072 6276 8084
rect 5951 8044 6276 8072
rect 5951 8041 5963 8044
rect 5905 8035 5963 8041
rect 6270 8032 6276 8044
rect 6328 8032 6334 8084
rect 3326 7896 3332 7948
rect 3384 7936 3390 7948
rect 4157 7939 4215 7945
rect 4157 7936 4169 7939
rect 3384 7908 4169 7936
rect 3384 7896 3390 7908
rect 4157 7905 4169 7908
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 1946 7828 1952 7880
rect 2004 7828 2010 7880
rect 2774 7760 2780 7812
rect 2832 7800 2838 7812
rect 3053 7803 3111 7809
rect 3053 7800 3065 7803
rect 2832 7772 3065 7800
rect 2832 7760 2838 7772
rect 3053 7769 3065 7772
rect 3099 7769 3111 7803
rect 3053 7763 3111 7769
rect 4430 7760 4436 7812
rect 4488 7760 4494 7812
rect 4982 7760 4988 7812
rect 5040 7760 5046 7812
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2682 7732 2688 7744
rect 1627 7704 2688 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 1104 7642 6670 7664
rect 1104 7590 2288 7642
rect 2340 7590 2352 7642
rect 2404 7590 2416 7642
rect 2468 7590 2480 7642
rect 2532 7590 2544 7642
rect 2596 7590 3644 7642
rect 3696 7590 3708 7642
rect 3760 7590 3772 7642
rect 3824 7590 3836 7642
rect 3888 7590 3900 7642
rect 3952 7590 5000 7642
rect 5052 7590 5064 7642
rect 5116 7590 5128 7642
rect 5180 7590 5192 7642
rect 5244 7590 5256 7642
rect 5308 7590 6356 7642
rect 6408 7590 6420 7642
rect 6472 7590 6484 7642
rect 6536 7590 6548 7642
rect 6600 7590 6612 7642
rect 6664 7590 6670 7642
rect 1104 7568 6670 7590
rect 1946 7528 1952 7540
rect 1780 7500 1952 7528
rect 1780 7378 1808 7500
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 3878 7488 3884 7540
rect 3936 7528 3942 7540
rect 4062 7528 4068 7540
rect 3936 7500 4068 7528
rect 3936 7488 3942 7500
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 4525 7531 4583 7537
rect 4525 7528 4537 7531
rect 4488 7500 4537 7528
rect 4488 7488 4494 7500
rect 4525 7497 4537 7500
rect 4571 7497 4583 7531
rect 4525 7491 4583 7497
rect 4890 7488 4896 7540
rect 4948 7488 4954 7540
rect 6086 7488 6092 7540
rect 6144 7528 6150 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 6144 7500 6193 7528
rect 6144 7488 6150 7500
rect 6181 7497 6193 7500
rect 6227 7497 6239 7531
rect 6181 7491 6239 7497
rect 2590 7420 2596 7472
rect 2648 7460 2654 7472
rect 4246 7460 4252 7472
rect 2648 7432 3464 7460
rect 2648 7420 2654 7432
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 3326 7392 3332 7404
rect 3191 7364 3332 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 3436 7401 3464 7432
rect 3712 7432 4252 7460
rect 3712 7401 3740 7432
rect 4246 7420 4252 7432
rect 4304 7420 4310 7472
rect 4908 7460 4936 7488
rect 4908 7432 5120 7460
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7361 3479 7395
rect 3421 7355 3479 7361
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 3237 7327 3295 7333
rect 3237 7324 3249 7327
rect 2915 7296 3249 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 3237 7293 3249 7296
rect 3283 7293 3295 7327
rect 3436 7324 3464 7355
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 4890 7392 4896 7404
rect 4847 7364 4896 7392
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 4356 7324 4384 7355
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 5092 7336 5120 7432
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 3436 7296 4384 7324
rect 3237 7287 3295 7293
rect 5074 7284 5080 7336
rect 5132 7284 5138 7336
rect 3510 7216 3516 7268
rect 3568 7216 3574 7268
rect 3602 7216 3608 7268
rect 3660 7216 3666 7268
rect 4157 7259 4215 7265
rect 4157 7225 4169 7259
rect 4203 7225 4215 7259
rect 4157 7219 4215 7225
rect 4249 7259 4307 7265
rect 4249 7225 4261 7259
rect 4295 7256 4307 7259
rect 4617 7259 4675 7265
rect 4617 7256 4629 7259
rect 4295 7228 4629 7256
rect 4295 7225 4307 7228
rect 4249 7219 4307 7225
rect 4617 7225 4629 7228
rect 4663 7225 4675 7259
rect 4617 7219 4675 7225
rect 1397 7191 1455 7197
rect 1397 7157 1409 7191
rect 1443 7188 1455 7191
rect 2222 7188 2228 7200
rect 1443 7160 2228 7188
rect 1443 7157 1455 7160
rect 1397 7151 1455 7157
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 4172 7188 4200 7219
rect 4338 7188 4344 7200
rect 4172 7160 4344 7188
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 4798 7148 4804 7200
rect 4856 7188 4862 7200
rect 4985 7191 5043 7197
rect 4985 7188 4997 7191
rect 4856 7160 4997 7188
rect 4856 7148 4862 7160
rect 4985 7157 4997 7160
rect 5031 7157 5043 7191
rect 4985 7151 5043 7157
rect 1104 7098 6532 7120
rect 1104 7046 1628 7098
rect 1680 7046 1692 7098
rect 1744 7046 1756 7098
rect 1808 7046 1820 7098
rect 1872 7046 1884 7098
rect 1936 7046 2984 7098
rect 3036 7046 3048 7098
rect 3100 7046 3112 7098
rect 3164 7046 3176 7098
rect 3228 7046 3240 7098
rect 3292 7046 4340 7098
rect 4392 7046 4404 7098
rect 4456 7046 4468 7098
rect 4520 7046 4532 7098
rect 4584 7046 4596 7098
rect 4648 7046 5696 7098
rect 5748 7046 5760 7098
rect 5812 7046 5824 7098
rect 5876 7046 5888 7098
rect 5940 7046 5952 7098
rect 6004 7046 6532 7098
rect 1104 7024 6532 7046
rect 2593 6987 2651 6993
rect 2593 6953 2605 6987
rect 2639 6984 2651 6987
rect 2774 6984 2780 6996
rect 2639 6956 2780 6984
rect 2639 6953 2651 6956
rect 2593 6947 2651 6953
rect 2774 6944 2780 6956
rect 2832 6944 2838 6996
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 3237 6987 3295 6993
rect 3237 6984 3249 6987
rect 3200 6956 3249 6984
rect 3200 6944 3206 6956
rect 3237 6953 3249 6956
rect 3283 6953 3295 6987
rect 3237 6947 3295 6953
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 3660 6956 3801 6984
rect 3660 6944 3666 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 3789 6947 3847 6953
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4341 6987 4399 6993
rect 4341 6984 4353 6987
rect 4304 6956 4353 6984
rect 4304 6944 4310 6956
rect 4341 6953 4353 6956
rect 4387 6953 4399 6987
rect 4341 6947 4399 6953
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 5442 6984 5448 6996
rect 4571 6956 5448 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 3160 6916 3188 6944
rect 4540 6916 4568 6947
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 1964 6888 4568 6916
rect 1578 6740 1584 6792
rect 1636 6740 1642 6792
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 1964 6780 1992 6888
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6848 2559 6851
rect 2869 6851 2927 6857
rect 2869 6848 2881 6851
rect 2547 6820 2881 6848
rect 2547 6817 2559 6820
rect 2501 6811 2559 6817
rect 2869 6817 2881 6820
rect 2915 6817 2927 6851
rect 2869 6811 2927 6817
rect 2958 6808 2964 6860
rect 3016 6808 3022 6860
rect 3068 6820 3464 6848
rect 1903 6752 1992 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 2038 6740 2044 6792
rect 2096 6740 2102 6792
rect 2130 6740 2136 6792
rect 2188 6740 2194 6792
rect 2222 6740 2228 6792
rect 2280 6780 2286 6792
rect 3068 6789 3096 6820
rect 3436 6792 3464 6820
rect 3878 6808 3884 6860
rect 3936 6808 3942 6860
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6848 4215 6851
rect 4246 6848 4252 6860
rect 4203 6820 4252 6848
rect 4203 6817 4215 6820
rect 4157 6811 4215 6817
rect 2317 6783 2375 6789
rect 2317 6780 2329 6783
rect 2280 6752 2329 6780
rect 2280 6740 2286 6752
rect 2317 6749 2329 6752
rect 2363 6749 2375 6783
rect 2317 6743 2375 6749
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6780 2835 6783
rect 3053 6783 3111 6789
rect 2823 6752 2912 6780
rect 2823 6749 2835 6752
rect 2777 6743 2835 6749
rect 1949 6715 2007 6721
rect 1949 6681 1961 6715
rect 1995 6712 2007 6715
rect 2590 6712 2596 6724
rect 1995 6684 2596 6712
rect 1995 6681 2007 6684
rect 1949 6675 2007 6681
rect 2590 6672 2596 6684
rect 2648 6712 2654 6724
rect 2884 6712 2912 6752
rect 3053 6749 3065 6783
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 3234 6740 3240 6792
rect 3292 6740 3298 6792
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 2648 6684 2912 6712
rect 3344 6712 3372 6743
rect 3418 6740 3424 6792
rect 3476 6740 3482 6792
rect 3896 6780 3924 6808
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3896 6752 3985 6780
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 4080 6780 4108 6811
rect 4246 6808 4252 6820
rect 4304 6848 4310 6860
rect 4890 6848 4896 6860
rect 4304 6820 4896 6848
rect 4304 6808 4310 6820
rect 4890 6808 4896 6820
rect 4948 6848 4954 6860
rect 6089 6851 6147 6857
rect 4948 6820 5856 6848
rect 4948 6808 4954 6820
rect 4522 6780 4528 6792
rect 4080 6752 4528 6780
rect 3973 6743 4031 6749
rect 3988 6712 4016 6743
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4246 6712 4252 6724
rect 3344 6684 3464 6712
rect 3988 6684 4252 6712
rect 2648 6672 2654 6684
rect 2884 6656 2912 6684
rect 3436 6656 3464 6684
rect 4246 6672 4252 6684
rect 4304 6672 4310 6724
rect 4632 6712 4660 6743
rect 4706 6740 4712 6792
rect 4764 6740 4770 6792
rect 5074 6740 5080 6792
rect 5132 6740 5138 6792
rect 5828 6789 5856 6820
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6178 6848 6184 6860
rect 6135 6820 6184 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 4890 6712 4896 6724
rect 4632 6684 4896 6712
rect 4890 6672 4896 6684
rect 4948 6712 4954 6724
rect 5092 6712 5120 6740
rect 4948 6684 5120 6712
rect 4948 6672 4954 6684
rect 2866 6604 2872 6656
rect 2924 6604 2930 6656
rect 3418 6604 3424 6656
rect 3476 6604 3482 6656
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 4062 6644 4068 6656
rect 3651 6616 4068 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 1104 6554 6670 6576
rect 1104 6502 2288 6554
rect 2340 6502 2352 6554
rect 2404 6502 2416 6554
rect 2468 6502 2480 6554
rect 2532 6502 2544 6554
rect 2596 6502 3644 6554
rect 3696 6502 3708 6554
rect 3760 6502 3772 6554
rect 3824 6502 3836 6554
rect 3888 6502 3900 6554
rect 3952 6502 5000 6554
rect 5052 6502 5064 6554
rect 5116 6502 5128 6554
rect 5180 6502 5192 6554
rect 5244 6502 5256 6554
rect 5308 6502 6356 6554
rect 6408 6502 6420 6554
rect 6472 6502 6484 6554
rect 6536 6502 6548 6554
rect 6600 6502 6612 6554
rect 6664 6502 6670 6554
rect 1104 6480 6670 6502
rect 1578 6400 1584 6452
rect 1636 6400 1642 6452
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 4062 6440 4068 6452
rect 2096 6412 4068 6440
rect 2096 6400 2102 6412
rect 4062 6400 4068 6412
rect 4120 6440 4126 6452
rect 4890 6440 4896 6452
rect 4120 6412 4896 6440
rect 4120 6400 4126 6412
rect 4890 6400 4896 6412
rect 4948 6440 4954 6452
rect 5077 6443 5135 6449
rect 5077 6440 5089 6443
rect 4948 6412 5089 6440
rect 4948 6400 4954 6412
rect 5077 6409 5089 6412
rect 5123 6440 5135 6443
rect 5442 6440 5448 6452
rect 5123 6412 5448 6440
rect 5123 6409 5135 6412
rect 5077 6403 5135 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 1596 6372 1624 6400
rect 1596 6344 2636 6372
rect 2056 6316 2084 6344
rect 1394 6264 1400 6316
rect 1452 6264 1458 6316
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 2608 6313 2636 6344
rect 4706 6332 4712 6384
rect 4764 6372 4770 6384
rect 4982 6372 4988 6384
rect 4764 6344 4988 6372
rect 4764 6332 4770 6344
rect 4982 6332 4988 6344
rect 5040 6372 5046 6384
rect 5040 6344 5948 6372
rect 5040 6332 5046 6344
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 2608 6236 2636 6267
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2832 6276 3065 6304
rect 2832 6264 2838 6276
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3418 6264 3424 6316
rect 3476 6304 3482 6316
rect 5920 6313 5948 6344
rect 4893 6307 4951 6313
rect 4893 6304 4905 6307
rect 3476 6276 4905 6304
rect 3476 6264 3482 6276
rect 4893 6273 4905 6276
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 3436 6236 3464 6264
rect 2608 6208 3464 6236
rect 4522 6196 4528 6248
rect 4580 6196 4586 6248
rect 2590 6128 2596 6180
rect 2648 6128 2654 6180
rect 2777 6171 2835 6177
rect 2777 6137 2789 6171
rect 2823 6168 2835 6171
rect 3418 6168 3424 6180
rect 2823 6140 3424 6168
rect 2823 6137 2835 6140
rect 2777 6131 2835 6137
rect 3418 6128 3424 6140
rect 3476 6168 3482 6180
rect 4540 6168 4568 6196
rect 4706 6168 4712 6180
rect 3476 6140 4712 6168
rect 3476 6128 3482 6140
rect 4706 6128 4712 6140
rect 4764 6128 4770 6180
rect 2608 6100 2636 6128
rect 3142 6100 3148 6112
rect 2608 6072 3148 6100
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4341 6103 4399 6109
rect 4341 6100 4353 6103
rect 4212 6072 4353 6100
rect 4212 6060 4218 6072
rect 4341 6069 4353 6072
rect 4387 6069 4399 6103
rect 4341 6063 4399 6069
rect 6086 6060 6092 6112
rect 6144 6060 6150 6112
rect 1104 6010 6532 6032
rect 1104 5958 1628 6010
rect 1680 5958 1692 6010
rect 1744 5958 1756 6010
rect 1808 5958 1820 6010
rect 1872 5958 1884 6010
rect 1936 5958 2984 6010
rect 3036 5958 3048 6010
rect 3100 5958 3112 6010
rect 3164 5958 3176 6010
rect 3228 5958 3240 6010
rect 3292 5958 4340 6010
rect 4392 5958 4404 6010
rect 4456 5958 4468 6010
rect 4520 5958 4532 6010
rect 4584 5958 4596 6010
rect 4648 5958 5696 6010
rect 5748 5958 5760 6010
rect 5812 5958 5824 6010
rect 5876 5958 5888 6010
rect 5940 5958 5952 6010
rect 6004 5958 6532 6010
rect 1104 5936 6532 5958
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3568 5868 3801 5896
rect 3568 5856 3574 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 4157 5899 4215 5905
rect 4157 5896 4169 5899
rect 3789 5859 3847 5865
rect 3896 5868 4169 5896
rect 3896 5760 3924 5868
rect 4157 5865 4169 5868
rect 4203 5896 4215 5899
rect 4798 5896 4804 5908
rect 4203 5868 4804 5896
rect 4203 5865 4215 5868
rect 4157 5859 4215 5865
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 4982 5856 4988 5908
rect 5040 5896 5046 5908
rect 5040 5868 5212 5896
rect 5040 5856 5046 5868
rect 4062 5788 4068 5840
rect 4120 5788 4126 5840
rect 4246 5788 4252 5840
rect 4304 5788 4310 5840
rect 4706 5788 4712 5840
rect 4764 5828 4770 5840
rect 4764 5800 5028 5828
rect 4764 5788 4770 5800
rect 3528 5732 3924 5760
rect 3528 5704 3556 5732
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 3510 5652 3516 5704
rect 3568 5652 3574 5704
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 4080 5692 4108 5788
rect 4264 5760 4292 5788
rect 4798 5760 4804 5772
rect 4264 5732 4804 5760
rect 4798 5720 4804 5732
rect 4856 5760 4862 5772
rect 5000 5769 5028 5800
rect 4893 5763 4951 5769
rect 4893 5760 4905 5763
rect 4856 5732 4905 5760
rect 4856 5720 4862 5732
rect 4893 5729 4905 5732
rect 4939 5729 4951 5763
rect 4893 5723 4951 5729
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5729 5043 5763
rect 4985 5723 5043 5729
rect 5095 5763 5153 5769
rect 5095 5729 5107 5763
rect 5141 5760 5153 5763
rect 5184 5760 5212 5868
rect 5141 5732 5212 5760
rect 5141 5729 5153 5732
rect 5095 5723 5153 5729
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 4080 5664 4261 5692
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 5813 5627 5871 5633
rect 5813 5593 5825 5627
rect 5859 5624 5871 5627
rect 6270 5624 6276 5636
rect 5859 5596 6276 5624
rect 5859 5593 5871 5596
rect 5813 5587 5871 5593
rect 6270 5584 6276 5596
rect 6328 5584 6334 5636
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 1946 5556 1952 5568
rect 1627 5528 1952 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 1946 5516 1952 5528
rect 2004 5516 2010 5568
rect 4706 5516 4712 5568
rect 4764 5516 4770 5568
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6178 5556 6184 5568
rect 6135 5528 6184 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 1104 5466 6670 5488
rect 1104 5414 2288 5466
rect 2340 5414 2352 5466
rect 2404 5414 2416 5466
rect 2468 5414 2480 5466
rect 2532 5414 2544 5466
rect 2596 5414 3644 5466
rect 3696 5414 3708 5466
rect 3760 5414 3772 5466
rect 3824 5414 3836 5466
rect 3888 5414 3900 5466
rect 3952 5414 5000 5466
rect 5052 5414 5064 5466
rect 5116 5414 5128 5466
rect 5180 5414 5192 5466
rect 5244 5414 5256 5466
rect 5308 5414 6356 5466
rect 6408 5414 6420 5466
rect 6472 5414 6484 5466
rect 6536 5414 6548 5466
rect 6600 5414 6612 5466
rect 6664 5414 6670 5466
rect 1104 5392 6670 5414
rect 2130 5352 2136 5364
rect 2056 5324 2136 5352
rect 2056 5293 2084 5324
rect 2130 5312 2136 5324
rect 2188 5352 2194 5364
rect 3510 5352 3516 5364
rect 2188 5324 3516 5352
rect 2188 5312 2194 5324
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 3804 5324 4200 5352
rect 2041 5287 2099 5293
rect 2041 5284 2053 5287
rect 1320 5256 2053 5284
rect 1320 5228 1348 5256
rect 2041 5253 2053 5256
rect 2087 5253 2099 5287
rect 2041 5247 2099 5253
rect 2498 5244 2504 5296
rect 2556 5284 2562 5296
rect 2866 5284 2872 5296
rect 2556 5256 2872 5284
rect 2556 5244 2562 5256
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 3804 5284 3832 5324
rect 4062 5284 4068 5296
rect 3160 5256 3832 5284
rect 3896 5256 4068 5284
rect 1302 5176 1308 5228
rect 1360 5176 1366 5228
rect 3160 5216 3188 5256
rect 2516 5188 3188 5216
rect 3237 5219 3295 5225
rect 2130 5108 2136 5160
rect 2188 5148 2194 5160
rect 2516 5157 2544 5188
rect 3237 5185 3249 5219
rect 3283 5216 3295 5219
rect 3326 5216 3332 5228
rect 3283 5188 3332 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 3418 5176 3424 5228
rect 3476 5176 3482 5228
rect 3510 5176 3516 5228
rect 3568 5176 3574 5228
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 2188 5120 2513 5148
rect 2188 5108 2194 5120
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 2590 5108 2596 5160
rect 2648 5108 2654 5160
rect 2961 5151 3019 5157
rect 2961 5117 2973 5151
rect 3007 5148 3019 5151
rect 3436 5148 3464 5176
rect 3896 5157 3924 5256
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 4172 5225 4200 5324
rect 4614 5312 4620 5364
rect 4672 5312 4678 5364
rect 4706 5312 4712 5364
rect 4764 5312 4770 5364
rect 4632 5225 4660 5312
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4629 5219 4687 5225
rect 4629 5185 4641 5219
rect 4675 5185 4687 5219
rect 4724 5216 4752 5312
rect 5534 5284 5540 5296
rect 4908 5256 5540 5284
rect 4908 5225 4936 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4724 5188 4813 5216
rect 4629 5179 4687 5185
rect 4801 5185 4813 5188
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5261 5219 5319 5225
rect 5040 5188 5212 5216
rect 5040 5176 5046 5188
rect 3007 5120 3464 5148
rect 3881 5151 3939 5157
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 3881 5117 3893 5151
rect 3927 5117 3939 5151
rect 3881 5111 3939 5117
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5148 4031 5151
rect 4246 5148 4252 5160
rect 4019 5120 4252 5148
rect 4019 5117 4031 5120
rect 3973 5111 4031 5117
rect 2038 5040 2044 5092
rect 2096 5040 2102 5092
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 3697 5083 3755 5089
rect 3697 5080 3709 5083
rect 3099 5052 3709 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 3697 5049 3709 5052
rect 3743 5080 3755 5083
rect 3988 5080 4016 5111
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 5077 5151 5135 5157
rect 5077 5148 5089 5151
rect 4755 5120 5089 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 5077 5117 5089 5120
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 4062 5080 4068 5092
rect 3743 5052 4068 5080
rect 3743 5049 3755 5052
rect 3697 5043 3755 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 4341 5083 4399 5089
rect 4341 5049 4353 5083
rect 4387 5080 4399 5083
rect 4798 5080 4804 5092
rect 4387 5052 4804 5080
rect 4387 5049 4399 5052
rect 4341 5043 4399 5049
rect 4798 5040 4804 5052
rect 4856 5040 4862 5092
rect 4982 5040 4988 5092
rect 5040 5040 5046 5092
rect 2682 4972 2688 5024
rect 2740 5012 2746 5024
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 2740 4984 2789 5012
rect 2740 4972 2746 4984
rect 2777 4981 2789 4984
rect 2823 4981 2835 5015
rect 2777 4975 2835 4981
rect 3418 4972 3424 5024
rect 3476 4972 3482 5024
rect 4433 5015 4491 5021
rect 4433 4981 4445 5015
rect 4479 5012 4491 5015
rect 5000 5012 5028 5040
rect 4479 4984 5028 5012
rect 5184 5012 5212 5188
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5307 5188 6009 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 5997 5185 6009 5188
rect 6043 5216 6055 5219
rect 6086 5216 6092 5228
rect 6043 5188 6092 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6086 5176 6092 5188
rect 6144 5176 6150 5228
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5500 5120 5549 5148
rect 5500 5108 5506 5120
rect 5537 5117 5549 5120
rect 5583 5148 5595 5151
rect 5905 5151 5963 5157
rect 5905 5148 5917 5151
rect 5583 5120 5917 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 5905 5117 5917 5120
rect 5951 5117 5963 5151
rect 5905 5111 5963 5117
rect 5350 5040 5356 5092
rect 5408 5080 5414 5092
rect 5629 5083 5687 5089
rect 5629 5080 5641 5083
rect 5408 5052 5641 5080
rect 5408 5040 5414 5052
rect 5629 5049 5641 5052
rect 5675 5049 5687 5083
rect 5629 5043 5687 5049
rect 5445 5015 5503 5021
rect 5445 5012 5457 5015
rect 5184 4984 5457 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 5445 4981 5457 4984
rect 5491 4981 5503 5015
rect 5445 4975 5503 4981
rect 5997 5015 6055 5021
rect 5997 4981 6009 5015
rect 6043 5012 6055 5015
rect 6362 5012 6368 5024
rect 6043 4984 6368 5012
rect 6043 4981 6055 4984
rect 5997 4975 6055 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 1104 4922 6532 4944
rect 1104 4870 1628 4922
rect 1680 4870 1692 4922
rect 1744 4870 1756 4922
rect 1808 4870 1820 4922
rect 1872 4870 1884 4922
rect 1936 4870 2984 4922
rect 3036 4870 3048 4922
rect 3100 4870 3112 4922
rect 3164 4870 3176 4922
rect 3228 4870 3240 4922
rect 3292 4870 4340 4922
rect 4392 4870 4404 4922
rect 4456 4870 4468 4922
rect 4520 4870 4532 4922
rect 4584 4870 4596 4922
rect 4648 4870 5696 4922
rect 5748 4870 5760 4922
rect 5812 4870 5824 4922
rect 5876 4870 5888 4922
rect 5940 4870 5952 4922
rect 6004 4870 6532 4922
rect 1104 4848 6532 4870
rect 3970 4808 3976 4820
rect 3896 4780 3976 4808
rect 2498 4700 2504 4752
rect 2556 4740 2562 4752
rect 2556 4712 3188 4740
rect 2556 4700 2562 4712
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 2516 4613 2544 4700
rect 2608 4613 2728 4638
rect 3160 4616 3188 4712
rect 3510 4632 3516 4684
rect 3568 4632 3574 4684
rect 3896 4681 3924 4780
rect 3970 4768 3976 4780
rect 4028 4808 4034 4820
rect 6270 4808 6276 4820
rect 4028 4780 6276 4808
rect 4028 4768 4034 4780
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 3881 4675 3939 4681
rect 3881 4641 3893 4675
rect 3927 4641 3939 4675
rect 3881 4635 3939 4641
rect 4062 4632 4068 4684
rect 4120 4632 4126 4684
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 4982 4672 4988 4684
rect 4663 4644 4988 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 2087 4607 2145 4613
rect 2087 4604 2099 4607
rect 2004 4576 2099 4604
rect 2004 4564 2010 4576
rect 2087 4573 2099 4576
rect 2133 4573 2145 4607
rect 2087 4567 2145 4573
rect 2472 4607 2544 4613
rect 2472 4573 2484 4607
rect 2518 4576 2544 4607
rect 2593 4610 2728 4613
rect 2593 4607 2651 4610
rect 2518 4573 2530 4576
rect 2472 4567 2530 4573
rect 2593 4573 2605 4607
rect 2639 4573 2651 4607
rect 2700 4604 2728 4610
rect 2958 4604 2964 4616
rect 2700 4576 2964 4604
rect 2593 4567 2651 4573
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 3142 4564 3148 4616
rect 3200 4564 3206 4616
rect 3234 4564 3240 4616
rect 3292 4564 3298 4616
rect 3528 4604 3556 4632
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3528 4576 3985 4604
rect 2225 4539 2283 4545
rect 2225 4505 2237 4539
rect 2271 4505 2283 4539
rect 2225 4499 2283 4505
rect 2317 4539 2375 4545
rect 2317 4505 2329 4539
rect 2363 4536 2375 4539
rect 2685 4539 2743 4545
rect 2685 4536 2697 4539
rect 2363 4508 2697 4536
rect 2363 4505 2375 4508
rect 2317 4499 2375 4505
rect 2685 4505 2697 4508
rect 2731 4505 2743 4539
rect 2685 4499 2743 4505
rect 1854 4428 1860 4480
rect 1912 4468 1918 4480
rect 1949 4471 2007 4477
rect 1949 4468 1961 4471
rect 1912 4440 1961 4468
rect 1912 4428 1918 4440
rect 1949 4437 1961 4440
rect 1995 4437 2007 4471
rect 2240 4468 2268 4499
rect 2866 4468 2872 4480
rect 2240 4440 2872 4468
rect 1949 4431 2007 4437
rect 2866 4428 2872 4440
rect 2924 4468 2930 4480
rect 3528 4468 3556 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 5258 4496 5264 4548
rect 5316 4496 5322 4548
rect 2924 4440 3556 4468
rect 2924 4428 2930 4440
rect 4246 4428 4252 4480
rect 4304 4428 4310 4480
rect 6089 4471 6147 4477
rect 6089 4437 6101 4471
rect 6135 4468 6147 4471
rect 6178 4468 6184 4480
rect 6135 4440 6184 4468
rect 6135 4437 6147 4440
rect 6089 4431 6147 4437
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 1104 4378 6670 4400
rect 1104 4326 2288 4378
rect 2340 4326 2352 4378
rect 2404 4326 2416 4378
rect 2468 4326 2480 4378
rect 2532 4326 2544 4378
rect 2596 4326 3644 4378
rect 3696 4326 3708 4378
rect 3760 4326 3772 4378
rect 3824 4326 3836 4378
rect 3888 4326 3900 4378
rect 3952 4326 5000 4378
rect 5052 4326 5064 4378
rect 5116 4326 5128 4378
rect 5180 4326 5192 4378
rect 5244 4326 5256 4378
rect 5308 4326 6356 4378
rect 6408 4326 6420 4378
rect 6472 4326 6484 4378
rect 6536 4326 6548 4378
rect 6600 4326 6612 4378
rect 6664 4326 6670 4378
rect 1104 4304 6670 4326
rect 3510 4224 3516 4276
rect 3568 4264 3574 4276
rect 4062 4264 4068 4276
rect 3568 4236 4068 4264
rect 3568 4224 3574 4236
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 3142 4156 3148 4208
rect 3200 4196 3206 4208
rect 4706 4196 4712 4208
rect 3200 4168 4712 4196
rect 3200 4156 3206 4168
rect 1486 4020 1492 4072
rect 1544 4020 1550 4072
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4060 1823 4063
rect 1854 4060 1860 4072
rect 1811 4032 1860 4060
rect 1811 4029 1823 4032
rect 1765 4023 1823 4029
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 2884 4060 2912 4114
rect 3418 4088 3424 4140
rect 3476 4088 3482 4140
rect 3528 4137 3556 4168
rect 3896 4140 3924 4168
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 4890 4156 4896 4208
rect 4948 4196 4954 4208
rect 4948 4168 5106 4196
rect 4948 4156 4954 4168
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 3789 4131 3847 4137
rect 3789 4128 3801 4131
rect 3752 4100 3801 4128
rect 3752 4088 3758 4100
rect 3789 4097 3801 4100
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 3878 4088 3884 4140
rect 3936 4088 3942 4140
rect 2958 4060 2964 4072
rect 2556 4032 2964 4060
rect 2556 4020 2562 4032
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3436 4060 3464 4088
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 3436 4032 3617 4060
rect 3605 4029 3617 4032
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 4338 4020 4344 4072
rect 4396 4020 4402 4072
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4060 4675 4063
rect 4706 4060 4712 4072
rect 4663 4032 4712 4060
rect 4663 4029 4675 4032
rect 4617 4023 4675 4029
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 3234 3952 3240 4004
rect 3292 3992 3298 4004
rect 3697 3995 3755 4001
rect 3292 3964 3464 3992
rect 3292 3952 3298 3964
rect 3326 3884 3332 3936
rect 3384 3884 3390 3936
rect 3436 3924 3464 3964
rect 3697 3961 3709 3995
rect 3743 3992 3755 3995
rect 3970 3992 3976 4004
rect 3743 3964 3976 3992
rect 3743 3961 3755 3964
rect 3697 3955 3755 3961
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 4062 3924 4068 3936
rect 3436 3896 4068 3924
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4356 3924 4384 4020
rect 5074 3924 5080 3936
rect 4356 3896 5080 3924
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 6086 3884 6092 3936
rect 6144 3884 6150 3936
rect 1104 3834 6532 3856
rect 1104 3782 1628 3834
rect 1680 3782 1692 3834
rect 1744 3782 1756 3834
rect 1808 3782 1820 3834
rect 1872 3782 1884 3834
rect 1936 3782 2984 3834
rect 3036 3782 3048 3834
rect 3100 3782 3112 3834
rect 3164 3782 3176 3834
rect 3228 3782 3240 3834
rect 3292 3782 4340 3834
rect 4392 3782 4404 3834
rect 4456 3782 4468 3834
rect 4520 3782 4532 3834
rect 4584 3782 4596 3834
rect 4648 3782 5696 3834
rect 5748 3782 5760 3834
rect 5812 3782 5824 3834
rect 5876 3782 5888 3834
rect 5940 3782 5952 3834
rect 6004 3782 6532 3834
rect 1104 3760 6532 3782
rect 1486 3680 1492 3732
rect 1544 3720 1550 3732
rect 1544 3692 3372 3720
rect 1544 3680 1550 3692
rect 3344 3593 3372 3692
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 4522 3720 4528 3732
rect 3936 3692 4528 3720
rect 3936 3680 3942 3692
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5074 3680 5080 3732
rect 5132 3680 5138 3732
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 5592 3692 5641 3720
rect 5592 3680 5598 3692
rect 5629 3689 5641 3692
rect 5675 3689 5687 3723
rect 5629 3683 5687 3689
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 6270 3720 6276 3732
rect 5868 3692 6276 3720
rect 5868 3680 5874 3692
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 3329 3587 3387 3593
rect 3329 3553 3341 3587
rect 3375 3584 3387 3587
rect 5092 3584 5120 3680
rect 3375 3556 5120 3584
rect 3375 3553 3387 3556
rect 3329 3547 3387 3553
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5500 3556 5917 3584
rect 5500 3544 5506 3556
rect 5905 3553 5917 3556
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 4154 3516 4160 3528
rect 3835 3488 4160 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 2498 3408 2504 3460
rect 2556 3408 2562 3460
rect 3053 3451 3111 3457
rect 3053 3417 3065 3451
rect 3099 3448 3111 3451
rect 3326 3448 3332 3460
rect 3099 3420 3332 3448
rect 3099 3417 3111 3420
rect 3053 3411 3111 3417
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 1578 3340 1584 3392
rect 1636 3340 1642 3392
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 5460 3380 5488 3544
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3516 6055 3519
rect 6178 3516 6184 3528
rect 6043 3488 6184 3516
rect 6043 3485 6055 3488
rect 5997 3479 6055 3485
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 3292 3352 5488 3380
rect 3292 3340 3298 3352
rect 1104 3290 6670 3312
rect 1104 3238 2288 3290
rect 2340 3238 2352 3290
rect 2404 3238 2416 3290
rect 2468 3238 2480 3290
rect 2532 3238 2544 3290
rect 2596 3238 3644 3290
rect 3696 3238 3708 3290
rect 3760 3238 3772 3290
rect 3824 3238 3836 3290
rect 3888 3238 3900 3290
rect 3952 3238 5000 3290
rect 5052 3238 5064 3290
rect 5116 3238 5128 3290
rect 5180 3238 5192 3290
rect 5244 3238 5256 3290
rect 5308 3238 6356 3290
rect 6408 3238 6420 3290
rect 6472 3238 6484 3290
rect 6536 3238 6548 3290
rect 6600 3238 6612 3290
rect 6664 3238 6670 3290
rect 1104 3216 6670 3238
rect 2866 3136 2872 3188
rect 2924 3136 2930 3188
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 3510 3176 3516 3188
rect 3467 3148 3516 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 3970 3176 3976 3188
rect 3835 3148 3976 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4706 3176 4712 3188
rect 4387 3148 4712 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 6089 3179 6147 3185
rect 6089 3145 6101 3179
rect 6135 3176 6147 3179
rect 6730 3176 6736 3188
rect 6135 3148 6736 3176
rect 6135 3145 6147 3148
rect 6089 3139 6147 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 2884 3108 2912 3136
rect 2884 3080 4108 3108
rect 934 3000 940 3052
rect 992 3040 998 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 992 3012 1409 3040
rect 992 3000 998 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 2130 3040 2136 3052
rect 1636 3012 2136 3040
rect 1636 3000 1642 3012
rect 2130 3000 2136 3012
rect 2188 3040 2194 3052
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2188 3012 3065 3040
rect 2188 3000 2194 3012
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 1673 2975 1731 2981
rect 1673 2972 1685 2975
rect 1360 2944 1685 2972
rect 1360 2932 1366 2944
rect 1673 2941 1685 2944
rect 1719 2941 1731 2975
rect 3068 2972 3096 3003
rect 3234 3000 3240 3052
rect 3292 3000 3298 3052
rect 3418 3000 3424 3052
rect 3476 3040 3482 3052
rect 4080 3049 4108 3080
rect 4172 3080 5948 3108
rect 4172 3049 4200 3080
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3476 3012 3985 3040
rect 3476 3000 3482 3012
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4246 3000 4252 3052
rect 4304 3000 4310 3052
rect 4522 3000 4528 3052
rect 4580 3000 4586 3052
rect 4837 3043 4895 3049
rect 4837 3009 4849 3043
rect 4883 3040 4895 3043
rect 5350 3040 5356 3052
rect 4883 3012 5356 3040
rect 4883 3009 4895 3012
rect 4837 3003 4895 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5920 3049 5948 3080
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 6086 3040 6092 3052
rect 5951 3012 6092 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 3326 2972 3332 2984
rect 3068 2944 3332 2972
rect 1673 2935 1731 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 4264 2972 4292 3000
rect 4709 2975 4767 2981
rect 4709 2972 4721 2975
rect 4264 2944 4721 2972
rect 4709 2941 4721 2944
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 4617 2907 4675 2913
rect 4617 2873 4629 2907
rect 4663 2904 4675 2907
rect 4798 2904 4804 2916
rect 4663 2876 4804 2904
rect 4663 2873 4675 2876
rect 4617 2867 4675 2873
rect 4798 2864 4804 2876
rect 4856 2864 4862 2916
rect 2682 2796 2688 2848
rect 2740 2836 2746 2848
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2740 2808 3065 2836
rect 2740 2796 2746 2808
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 3053 2799 3111 2805
rect 1104 2746 6532 2768
rect 1104 2694 1628 2746
rect 1680 2694 1692 2746
rect 1744 2694 1756 2746
rect 1808 2694 1820 2746
rect 1872 2694 1884 2746
rect 1936 2694 2984 2746
rect 3036 2694 3048 2746
rect 3100 2694 3112 2746
rect 3164 2694 3176 2746
rect 3228 2694 3240 2746
rect 3292 2694 4340 2746
rect 4392 2694 4404 2746
rect 4456 2694 4468 2746
rect 4520 2694 4532 2746
rect 4584 2694 4596 2746
rect 4648 2694 5696 2746
rect 5748 2694 5760 2746
rect 5812 2694 5824 2746
rect 5876 2694 5888 2746
rect 5940 2694 5952 2746
rect 6004 2694 6532 2746
rect 1104 2672 6532 2694
rect 3326 2388 3332 2440
rect 3384 2428 3390 2440
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 3384 2400 5365 2428
rect 3384 2388 3390 2400
rect 5353 2397 5365 2400
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 4062 2320 4068 2372
rect 4120 2360 4126 2372
rect 5813 2363 5871 2369
rect 5813 2360 5825 2363
rect 4120 2332 5825 2360
rect 4120 2320 4126 2332
rect 5813 2329 5825 2332
rect 5859 2329 5871 2363
rect 5813 2323 5871 2329
rect 5534 2252 5540 2304
rect 5592 2252 5598 2304
rect 6089 2295 6147 2301
rect 6089 2261 6101 2295
rect 6135 2292 6147 2295
rect 6178 2292 6184 2304
rect 6135 2264 6184 2292
rect 6135 2261 6147 2264
rect 6089 2255 6147 2261
rect 6178 2252 6184 2264
rect 6236 2252 6242 2304
rect 1104 2202 6670 2224
rect 1104 2150 2288 2202
rect 2340 2150 2352 2202
rect 2404 2150 2416 2202
rect 2468 2150 2480 2202
rect 2532 2150 2544 2202
rect 2596 2150 3644 2202
rect 3696 2150 3708 2202
rect 3760 2150 3772 2202
rect 3824 2150 3836 2202
rect 3888 2150 3900 2202
rect 3952 2150 5000 2202
rect 5052 2150 5064 2202
rect 5116 2150 5128 2202
rect 5180 2150 5192 2202
rect 5244 2150 5256 2202
rect 5308 2150 6356 2202
rect 6408 2150 6420 2202
rect 6472 2150 6484 2202
rect 6536 2150 6548 2202
rect 6600 2150 6612 2202
rect 6664 2150 6670 2202
rect 1104 2128 6670 2150
<< via1 >>
rect 1628 10310 1680 10362
rect 1692 10310 1744 10362
rect 1756 10310 1808 10362
rect 1820 10310 1872 10362
rect 1884 10310 1936 10362
rect 2984 10310 3036 10362
rect 3048 10310 3100 10362
rect 3112 10310 3164 10362
rect 3176 10310 3228 10362
rect 3240 10310 3292 10362
rect 4340 10310 4392 10362
rect 4404 10310 4456 10362
rect 4468 10310 4520 10362
rect 4532 10310 4584 10362
rect 4596 10310 4648 10362
rect 5696 10310 5748 10362
rect 5760 10310 5812 10362
rect 5824 10310 5876 10362
rect 5888 10310 5940 10362
rect 5952 10310 6004 10362
rect 5356 10251 5408 10260
rect 5356 10217 5365 10251
rect 5365 10217 5399 10251
rect 5399 10217 5408 10251
rect 5356 10208 5408 10217
rect 6368 10208 6420 10260
rect 940 10004 992 10056
rect 5448 10004 5500 10056
rect 5356 9936 5408 9988
rect 3516 9868 3568 9920
rect 2288 9766 2340 9818
rect 2352 9766 2404 9818
rect 2416 9766 2468 9818
rect 2480 9766 2532 9818
rect 2544 9766 2596 9818
rect 3644 9766 3696 9818
rect 3708 9766 3760 9818
rect 3772 9766 3824 9818
rect 3836 9766 3888 9818
rect 3900 9766 3952 9818
rect 5000 9766 5052 9818
rect 5064 9766 5116 9818
rect 5128 9766 5180 9818
rect 5192 9766 5244 9818
rect 5256 9766 5308 9818
rect 6356 9766 6408 9818
rect 6420 9766 6472 9818
rect 6484 9766 6536 9818
rect 6548 9766 6600 9818
rect 6612 9766 6664 9818
rect 5356 9707 5408 9716
rect 5356 9673 5365 9707
rect 5365 9673 5399 9707
rect 5399 9673 5408 9707
rect 5356 9664 5408 9673
rect 4252 9596 4304 9648
rect 940 9528 992 9580
rect 2688 9528 2740 9580
rect 4896 9460 4948 9512
rect 5356 9460 5408 9512
rect 6092 9596 6144 9648
rect 6276 9528 6328 9580
rect 6184 9392 6236 9444
rect 1952 9324 2004 9376
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 3516 9324 3568 9376
rect 5448 9324 5500 9376
rect 6736 9324 6788 9376
rect 1628 9222 1680 9274
rect 1692 9222 1744 9274
rect 1756 9222 1808 9274
rect 1820 9222 1872 9274
rect 1884 9222 1936 9274
rect 2984 9222 3036 9274
rect 3048 9222 3100 9274
rect 3112 9222 3164 9274
rect 3176 9222 3228 9274
rect 3240 9222 3292 9274
rect 4340 9222 4392 9274
rect 4404 9222 4456 9274
rect 4468 9222 4520 9274
rect 4532 9222 4584 9274
rect 4596 9222 4648 9274
rect 5696 9222 5748 9274
rect 5760 9222 5812 9274
rect 5824 9222 5876 9274
rect 5888 9222 5940 9274
rect 5952 9222 6004 9274
rect 5448 9120 5500 9172
rect 4252 9052 4304 9104
rect 6092 9052 6144 9104
rect 6184 9052 6236 9104
rect 3516 8959 3568 8968
rect 3516 8925 3525 8959
rect 3525 8925 3559 8959
rect 3559 8925 3568 8959
rect 3516 8916 3568 8925
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4712 8984 4764 9036
rect 5356 8848 5408 8900
rect 6092 8916 6144 8968
rect 2872 8780 2924 8832
rect 4252 8780 4304 8832
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 2288 8678 2340 8730
rect 2352 8678 2404 8730
rect 2416 8678 2468 8730
rect 2480 8678 2532 8730
rect 2544 8678 2596 8730
rect 3644 8678 3696 8730
rect 3708 8678 3760 8730
rect 3772 8678 3824 8730
rect 3836 8678 3888 8730
rect 3900 8678 3952 8730
rect 5000 8678 5052 8730
rect 5064 8678 5116 8730
rect 5128 8678 5180 8730
rect 5192 8678 5244 8730
rect 5256 8678 5308 8730
rect 6356 8678 6408 8730
rect 6420 8678 6472 8730
rect 6484 8678 6536 8730
rect 6548 8678 6600 8730
rect 6612 8678 6664 8730
rect 1952 8508 2004 8560
rect 4988 8508 5040 8560
rect 4160 8440 4212 8492
rect 4804 8372 4856 8424
rect 3332 8236 3384 8288
rect 1628 8134 1680 8186
rect 1692 8134 1744 8186
rect 1756 8134 1808 8186
rect 1820 8134 1872 8186
rect 1884 8134 1936 8186
rect 2984 8134 3036 8186
rect 3048 8134 3100 8186
rect 3112 8134 3164 8186
rect 3176 8134 3228 8186
rect 3240 8134 3292 8186
rect 4340 8134 4392 8186
rect 4404 8134 4456 8186
rect 4468 8134 4520 8186
rect 4532 8134 4584 8186
rect 4596 8134 4648 8186
rect 5696 8134 5748 8186
rect 5760 8134 5812 8186
rect 5824 8134 5876 8186
rect 5888 8134 5940 8186
rect 5952 8134 6004 8186
rect 3240 8032 3292 8084
rect 3516 8032 3568 8084
rect 5632 8032 5684 8084
rect 6276 8032 6328 8084
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 1952 7828 2004 7880
rect 2780 7760 2832 7812
rect 4436 7803 4488 7812
rect 4436 7769 4445 7803
rect 4445 7769 4479 7803
rect 4479 7769 4488 7803
rect 4436 7760 4488 7769
rect 4988 7760 5040 7812
rect 2688 7692 2740 7744
rect 2288 7590 2340 7642
rect 2352 7590 2404 7642
rect 2416 7590 2468 7642
rect 2480 7590 2532 7642
rect 2544 7590 2596 7642
rect 3644 7590 3696 7642
rect 3708 7590 3760 7642
rect 3772 7590 3824 7642
rect 3836 7590 3888 7642
rect 3900 7590 3952 7642
rect 5000 7590 5052 7642
rect 5064 7590 5116 7642
rect 5128 7590 5180 7642
rect 5192 7590 5244 7642
rect 5256 7590 5308 7642
rect 6356 7590 6408 7642
rect 6420 7590 6472 7642
rect 6484 7590 6536 7642
rect 6548 7590 6600 7642
rect 6612 7590 6664 7642
rect 1952 7488 2004 7540
rect 3884 7488 3936 7540
rect 4068 7488 4120 7540
rect 4436 7488 4488 7540
rect 4896 7488 4948 7540
rect 6092 7488 6144 7540
rect 2596 7420 2648 7472
rect 3332 7352 3384 7404
rect 4252 7420 4304 7472
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 4896 7352 4948 7404
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 5080 7327 5132 7336
rect 5080 7293 5089 7327
rect 5089 7293 5123 7327
rect 5123 7293 5132 7327
rect 5080 7284 5132 7293
rect 3516 7259 3568 7268
rect 3516 7225 3525 7259
rect 3525 7225 3559 7259
rect 3559 7225 3568 7259
rect 3516 7216 3568 7225
rect 3608 7259 3660 7268
rect 3608 7225 3617 7259
rect 3617 7225 3651 7259
rect 3651 7225 3660 7259
rect 3608 7216 3660 7225
rect 2228 7148 2280 7200
rect 4344 7148 4396 7200
rect 4804 7148 4856 7200
rect 1628 7046 1680 7098
rect 1692 7046 1744 7098
rect 1756 7046 1808 7098
rect 1820 7046 1872 7098
rect 1884 7046 1936 7098
rect 2984 7046 3036 7098
rect 3048 7046 3100 7098
rect 3112 7046 3164 7098
rect 3176 7046 3228 7098
rect 3240 7046 3292 7098
rect 4340 7046 4392 7098
rect 4404 7046 4456 7098
rect 4468 7046 4520 7098
rect 4532 7046 4584 7098
rect 4596 7046 4648 7098
rect 5696 7046 5748 7098
rect 5760 7046 5812 7098
rect 5824 7046 5876 7098
rect 5888 7046 5940 7098
rect 5952 7046 6004 7098
rect 2780 6944 2832 6996
rect 3148 6944 3200 6996
rect 3608 6944 3660 6996
rect 4252 6944 4304 6996
rect 5448 6944 5500 6996
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 2964 6851 3016 6860
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 2964 6808 3016 6817
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 2228 6740 2280 6792
rect 3884 6808 3936 6860
rect 2596 6672 2648 6724
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 3424 6740 3476 6792
rect 4252 6808 4304 6860
rect 4896 6808 4948 6860
rect 4528 6740 4580 6792
rect 4252 6672 4304 6724
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 5080 6740 5132 6792
rect 6184 6808 6236 6860
rect 4896 6672 4948 6724
rect 2872 6604 2924 6656
rect 3424 6604 3476 6656
rect 4068 6604 4120 6656
rect 2288 6502 2340 6554
rect 2352 6502 2404 6554
rect 2416 6502 2468 6554
rect 2480 6502 2532 6554
rect 2544 6502 2596 6554
rect 3644 6502 3696 6554
rect 3708 6502 3760 6554
rect 3772 6502 3824 6554
rect 3836 6502 3888 6554
rect 3900 6502 3952 6554
rect 5000 6502 5052 6554
rect 5064 6502 5116 6554
rect 5128 6502 5180 6554
rect 5192 6502 5244 6554
rect 5256 6502 5308 6554
rect 6356 6502 6408 6554
rect 6420 6502 6472 6554
rect 6484 6502 6536 6554
rect 6548 6502 6600 6554
rect 6612 6502 6664 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2044 6400 2096 6452
rect 4068 6400 4120 6452
rect 4896 6400 4948 6452
rect 5448 6400 5500 6452
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 2044 6264 2096 6316
rect 4712 6332 4764 6384
rect 4988 6332 5040 6384
rect 2780 6264 2832 6316
rect 3424 6264 3476 6316
rect 4528 6196 4580 6248
rect 2596 6128 2648 6180
rect 3424 6128 3476 6180
rect 4712 6128 4764 6180
rect 3148 6060 3200 6112
rect 4160 6060 4212 6112
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 1628 5958 1680 6010
rect 1692 5958 1744 6010
rect 1756 5958 1808 6010
rect 1820 5958 1872 6010
rect 1884 5958 1936 6010
rect 2984 5958 3036 6010
rect 3048 5958 3100 6010
rect 3112 5958 3164 6010
rect 3176 5958 3228 6010
rect 3240 5958 3292 6010
rect 4340 5958 4392 6010
rect 4404 5958 4456 6010
rect 4468 5958 4520 6010
rect 4532 5958 4584 6010
rect 4596 5958 4648 6010
rect 5696 5958 5748 6010
rect 5760 5958 5812 6010
rect 5824 5958 5876 6010
rect 5888 5958 5940 6010
rect 5952 5958 6004 6010
rect 3516 5856 3568 5908
rect 4804 5856 4856 5908
rect 4988 5856 5040 5908
rect 4068 5788 4120 5840
rect 4252 5788 4304 5840
rect 4712 5788 4764 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 3516 5652 3568 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 4804 5720 4856 5772
rect 6276 5584 6328 5636
rect 1952 5516 2004 5568
rect 4712 5559 4764 5568
rect 4712 5525 4721 5559
rect 4721 5525 4755 5559
rect 4755 5525 4764 5559
rect 4712 5516 4764 5525
rect 6184 5516 6236 5568
rect 2288 5414 2340 5466
rect 2352 5414 2404 5466
rect 2416 5414 2468 5466
rect 2480 5414 2532 5466
rect 2544 5414 2596 5466
rect 3644 5414 3696 5466
rect 3708 5414 3760 5466
rect 3772 5414 3824 5466
rect 3836 5414 3888 5466
rect 3900 5414 3952 5466
rect 5000 5414 5052 5466
rect 5064 5414 5116 5466
rect 5128 5414 5180 5466
rect 5192 5414 5244 5466
rect 5256 5414 5308 5466
rect 6356 5414 6408 5466
rect 6420 5414 6472 5466
rect 6484 5414 6536 5466
rect 6548 5414 6600 5466
rect 6612 5414 6664 5466
rect 2136 5312 2188 5364
rect 3516 5312 3568 5364
rect 2504 5244 2556 5296
rect 2872 5244 2924 5296
rect 1308 5176 1360 5228
rect 2136 5108 2188 5160
rect 3332 5176 3384 5228
rect 3424 5176 3476 5228
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 2596 5151 2648 5160
rect 2596 5117 2605 5151
rect 2605 5117 2639 5151
rect 2639 5117 2648 5151
rect 2596 5108 2648 5117
rect 4068 5244 4120 5296
rect 4620 5312 4672 5364
rect 4712 5312 4764 5364
rect 5540 5244 5592 5296
rect 4988 5176 5040 5228
rect 2044 5083 2096 5092
rect 2044 5049 2053 5083
rect 2053 5049 2087 5083
rect 2087 5049 2096 5083
rect 2044 5040 2096 5049
rect 4252 5108 4304 5160
rect 4068 5040 4120 5092
rect 4804 5040 4856 5092
rect 4988 5040 5040 5092
rect 2688 4972 2740 5024
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 6092 5176 6144 5228
rect 5448 5108 5500 5160
rect 5356 5040 5408 5092
rect 6368 4972 6420 5024
rect 1628 4870 1680 4922
rect 1692 4870 1744 4922
rect 1756 4870 1808 4922
rect 1820 4870 1872 4922
rect 1884 4870 1936 4922
rect 2984 4870 3036 4922
rect 3048 4870 3100 4922
rect 3112 4870 3164 4922
rect 3176 4870 3228 4922
rect 3240 4870 3292 4922
rect 4340 4870 4392 4922
rect 4404 4870 4456 4922
rect 4468 4870 4520 4922
rect 4532 4870 4584 4922
rect 4596 4870 4648 4922
rect 5696 4870 5748 4922
rect 5760 4870 5812 4922
rect 5824 4870 5876 4922
rect 5888 4870 5940 4922
rect 5952 4870 6004 4922
rect 2504 4700 2556 4752
rect 1952 4564 2004 4616
rect 3516 4632 3568 4684
rect 3976 4768 4028 4820
rect 6276 4768 6328 4820
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 4988 4632 5040 4684
rect 2964 4564 3016 4616
rect 3148 4564 3200 4616
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 1860 4428 1912 4480
rect 2872 4428 2924 4480
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 5264 4496 5316 4548
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 6184 4428 6236 4480
rect 2288 4326 2340 4378
rect 2352 4326 2404 4378
rect 2416 4326 2468 4378
rect 2480 4326 2532 4378
rect 2544 4326 2596 4378
rect 3644 4326 3696 4378
rect 3708 4326 3760 4378
rect 3772 4326 3824 4378
rect 3836 4326 3888 4378
rect 3900 4326 3952 4378
rect 5000 4326 5052 4378
rect 5064 4326 5116 4378
rect 5128 4326 5180 4378
rect 5192 4326 5244 4378
rect 5256 4326 5308 4378
rect 6356 4326 6408 4378
rect 6420 4326 6472 4378
rect 6484 4326 6536 4378
rect 6548 4326 6600 4378
rect 6612 4326 6664 4378
rect 3516 4224 3568 4276
rect 4068 4224 4120 4276
rect 3148 4156 3200 4208
rect 1492 4063 1544 4072
rect 1492 4029 1501 4063
rect 1501 4029 1535 4063
rect 1535 4029 1544 4063
rect 1492 4020 1544 4029
rect 1860 4020 1912 4072
rect 2504 4020 2556 4072
rect 3424 4088 3476 4140
rect 4712 4156 4764 4208
rect 4896 4156 4948 4208
rect 3700 4088 3752 4140
rect 3884 4088 3936 4140
rect 2964 4020 3016 4072
rect 4344 4063 4396 4072
rect 4344 4029 4353 4063
rect 4353 4029 4387 4063
rect 4387 4029 4396 4063
rect 4344 4020 4396 4029
rect 4712 4020 4764 4072
rect 3240 3995 3292 4004
rect 3240 3961 3249 3995
rect 3249 3961 3283 3995
rect 3283 3961 3292 3995
rect 3240 3952 3292 3961
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 3332 3884 3384 3893
rect 3976 3952 4028 4004
rect 4068 3884 4120 3936
rect 5080 3884 5132 3936
rect 6092 3927 6144 3936
rect 6092 3893 6101 3927
rect 6101 3893 6135 3927
rect 6135 3893 6144 3927
rect 6092 3884 6144 3893
rect 1628 3782 1680 3834
rect 1692 3782 1744 3834
rect 1756 3782 1808 3834
rect 1820 3782 1872 3834
rect 1884 3782 1936 3834
rect 2984 3782 3036 3834
rect 3048 3782 3100 3834
rect 3112 3782 3164 3834
rect 3176 3782 3228 3834
rect 3240 3782 3292 3834
rect 4340 3782 4392 3834
rect 4404 3782 4456 3834
rect 4468 3782 4520 3834
rect 4532 3782 4584 3834
rect 4596 3782 4648 3834
rect 5696 3782 5748 3834
rect 5760 3782 5812 3834
rect 5824 3782 5876 3834
rect 5888 3782 5940 3834
rect 5952 3782 6004 3834
rect 1492 3680 1544 3732
rect 3884 3680 3936 3732
rect 4528 3680 4580 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 5540 3680 5592 3732
rect 5816 3723 5868 3732
rect 5816 3689 5825 3723
rect 5825 3689 5859 3723
rect 5859 3689 5868 3723
rect 5816 3680 5868 3689
rect 6276 3680 6328 3732
rect 5448 3544 5500 3596
rect 4160 3476 4212 3528
rect 2504 3408 2556 3460
rect 3332 3408 3384 3460
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 3240 3340 3292 3392
rect 6184 3476 6236 3528
rect 2288 3238 2340 3290
rect 2352 3238 2404 3290
rect 2416 3238 2468 3290
rect 2480 3238 2532 3290
rect 2544 3238 2596 3290
rect 3644 3238 3696 3290
rect 3708 3238 3760 3290
rect 3772 3238 3824 3290
rect 3836 3238 3888 3290
rect 3900 3238 3952 3290
rect 5000 3238 5052 3290
rect 5064 3238 5116 3290
rect 5128 3238 5180 3290
rect 5192 3238 5244 3290
rect 5256 3238 5308 3290
rect 6356 3238 6408 3290
rect 6420 3238 6472 3290
rect 6484 3238 6536 3290
rect 6548 3238 6600 3290
rect 6612 3238 6664 3290
rect 2872 3136 2924 3188
rect 3516 3136 3568 3188
rect 3976 3136 4028 3188
rect 4712 3136 4764 3188
rect 6736 3136 6788 3188
rect 940 3000 992 3052
rect 1584 3000 1636 3052
rect 2136 3000 2188 3052
rect 1308 2932 1360 2984
rect 3240 3043 3292 3052
rect 3240 3009 3249 3043
rect 3249 3009 3283 3043
rect 3283 3009 3292 3043
rect 3240 3000 3292 3009
rect 3424 3000 3476 3052
rect 4252 3000 4304 3052
rect 4528 3043 4580 3052
rect 4528 3009 4537 3043
rect 4537 3009 4571 3043
rect 4571 3009 4580 3043
rect 4528 3000 4580 3009
rect 5356 3000 5408 3052
rect 6092 3000 6144 3052
rect 3332 2932 3384 2984
rect 4804 2864 4856 2916
rect 2688 2796 2740 2848
rect 1628 2694 1680 2746
rect 1692 2694 1744 2746
rect 1756 2694 1808 2746
rect 1820 2694 1872 2746
rect 1884 2694 1936 2746
rect 2984 2694 3036 2746
rect 3048 2694 3100 2746
rect 3112 2694 3164 2746
rect 3176 2694 3228 2746
rect 3240 2694 3292 2746
rect 4340 2694 4392 2746
rect 4404 2694 4456 2746
rect 4468 2694 4520 2746
rect 4532 2694 4584 2746
rect 4596 2694 4648 2746
rect 5696 2694 5748 2746
rect 5760 2694 5812 2746
rect 5824 2694 5876 2746
rect 5888 2694 5940 2746
rect 5952 2694 6004 2746
rect 3332 2388 3384 2440
rect 4068 2320 4120 2372
rect 5540 2295 5592 2304
rect 5540 2261 5549 2295
rect 5549 2261 5583 2295
rect 5583 2261 5592 2295
rect 5540 2252 5592 2261
rect 6184 2252 6236 2304
rect 2288 2150 2340 2202
rect 2352 2150 2404 2202
rect 2416 2150 2468 2202
rect 2480 2150 2532 2202
rect 2544 2150 2596 2202
rect 3644 2150 3696 2202
rect 3708 2150 3760 2202
rect 3772 2150 3824 2202
rect 3836 2150 3888 2202
rect 3900 2150 3952 2202
rect 5000 2150 5052 2202
rect 5064 2150 5116 2202
rect 5128 2150 5180 2202
rect 5192 2150 5244 2202
rect 5256 2150 5308 2202
rect 6356 2150 6408 2202
rect 6420 2150 6472 2202
rect 6484 2150 6536 2202
rect 6548 2150 6600 2202
rect 6612 2150 6664 2202
<< metal2 >>
rect 6366 11520 6422 11529
rect 6366 11455 6422 11464
rect 938 10976 994 10985
rect 938 10911 994 10920
rect 952 10062 980 10911
rect 1628 10364 1936 10373
rect 1628 10362 1634 10364
rect 1690 10362 1714 10364
rect 1770 10362 1794 10364
rect 1850 10362 1874 10364
rect 1930 10362 1936 10364
rect 1690 10310 1692 10362
rect 1872 10310 1874 10362
rect 1628 10308 1634 10310
rect 1690 10308 1714 10310
rect 1770 10308 1794 10310
rect 1850 10308 1874 10310
rect 1930 10308 1936 10310
rect 1628 10299 1936 10308
rect 2984 10364 3292 10373
rect 2984 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3150 10364
rect 3206 10362 3230 10364
rect 3286 10362 3292 10364
rect 3046 10310 3048 10362
rect 3228 10310 3230 10362
rect 2984 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3150 10310
rect 3206 10308 3230 10310
rect 3286 10308 3292 10310
rect 2984 10299 3292 10308
rect 4340 10364 4648 10373
rect 4340 10362 4346 10364
rect 4402 10362 4426 10364
rect 4482 10362 4506 10364
rect 4562 10362 4586 10364
rect 4642 10362 4648 10364
rect 4402 10310 4404 10362
rect 4584 10310 4586 10362
rect 4340 10308 4346 10310
rect 4402 10308 4426 10310
rect 4482 10308 4506 10310
rect 4562 10308 4586 10310
rect 4642 10308 4648 10310
rect 4340 10299 4648 10308
rect 5696 10364 6004 10373
rect 5696 10362 5702 10364
rect 5758 10362 5782 10364
rect 5838 10362 5862 10364
rect 5918 10362 5942 10364
rect 5998 10362 6004 10364
rect 5758 10310 5760 10362
rect 5940 10310 5942 10362
rect 5696 10308 5702 10310
rect 5758 10308 5782 10310
rect 5838 10308 5862 10310
rect 5918 10308 5942 10310
rect 5998 10308 6004 10310
rect 5696 10299 6004 10308
rect 6380 10266 6408 11455
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 5368 10169 5396 10202
rect 5354 10160 5410 10169
rect 5354 10095 5410 10104
rect 940 10056 992 10062
rect 940 9998 992 10004
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 2288 9820 2596 9829
rect 2288 9818 2294 9820
rect 2350 9818 2374 9820
rect 2430 9818 2454 9820
rect 2510 9818 2534 9820
rect 2590 9818 2596 9820
rect 2350 9766 2352 9818
rect 2532 9766 2534 9818
rect 2288 9764 2294 9766
rect 2350 9764 2374 9766
rect 2430 9764 2454 9766
rect 2510 9764 2534 9766
rect 2590 9764 2596 9766
rect 2288 9755 2596 9764
rect 940 9580 992 9586
rect 940 9522 992 9528
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 952 9081 980 9522
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1628 9276 1936 9285
rect 1628 9274 1634 9276
rect 1690 9274 1714 9276
rect 1770 9274 1794 9276
rect 1850 9274 1874 9276
rect 1930 9274 1936 9276
rect 1690 9222 1692 9274
rect 1872 9222 1874 9274
rect 1628 9220 1634 9222
rect 1690 9220 1714 9222
rect 1770 9220 1794 9222
rect 1850 9220 1874 9222
rect 1930 9220 1936 9222
rect 1628 9211 1936 9220
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 1964 8566 1992 9318
rect 2288 8732 2596 8741
rect 2288 8730 2294 8732
rect 2350 8730 2374 8732
rect 2430 8730 2454 8732
rect 2510 8730 2534 8732
rect 2590 8730 2596 8732
rect 2350 8678 2352 8730
rect 2532 8678 2534 8730
rect 2288 8676 2294 8678
rect 2350 8676 2374 8678
rect 2430 8676 2454 8678
rect 2510 8676 2534 8678
rect 2590 8676 2596 8678
rect 2288 8667 2596 8676
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 1628 8188 1936 8197
rect 1628 8186 1634 8188
rect 1690 8186 1714 8188
rect 1770 8186 1794 8188
rect 1850 8186 1874 8188
rect 1930 8186 1936 8188
rect 1690 8134 1692 8186
rect 1872 8134 1874 8186
rect 1628 8132 1634 8134
rect 1690 8132 1714 8134
rect 1770 8132 1794 8134
rect 1850 8132 1874 8134
rect 1930 8132 1936 8134
rect 1628 8123 1936 8132
rect 1964 7886 1992 8502
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1964 7546 1992 7822
rect 2700 7750 2728 9522
rect 3528 9382 3556 9862
rect 3644 9820 3952 9829
rect 3644 9818 3650 9820
rect 3706 9818 3730 9820
rect 3786 9818 3810 9820
rect 3866 9818 3890 9820
rect 3946 9818 3952 9820
rect 3706 9766 3708 9818
rect 3888 9766 3890 9818
rect 3644 9764 3650 9766
rect 3706 9764 3730 9766
rect 3786 9764 3810 9766
rect 3866 9764 3890 9766
rect 3946 9764 3952 9766
rect 3644 9755 3952 9764
rect 5000 9820 5308 9829
rect 5000 9818 5006 9820
rect 5062 9818 5086 9820
rect 5142 9818 5166 9820
rect 5222 9818 5246 9820
rect 5302 9818 5308 9820
rect 5062 9766 5064 9818
rect 5244 9766 5246 9818
rect 5000 9764 5006 9766
rect 5062 9764 5086 9766
rect 5142 9764 5166 9766
rect 5222 9764 5246 9766
rect 5302 9764 5308 9766
rect 5000 9755 5308 9764
rect 5368 9722 5396 9930
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 4252 9648 4304 9654
rect 5460 9602 5488 9998
rect 6356 9820 6664 9829
rect 6356 9818 6362 9820
rect 6418 9818 6442 9820
rect 6498 9818 6522 9820
rect 6578 9818 6602 9820
rect 6658 9818 6664 9820
rect 6418 9766 6420 9818
rect 6600 9766 6602 9818
rect 6356 9764 6362 9766
rect 6418 9764 6442 9766
rect 6498 9764 6522 9766
rect 6578 9764 6602 9766
rect 6658 9764 6664 9766
rect 6356 9755 6664 9764
rect 4252 9590 4304 9596
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 2984 9276 3292 9285
rect 2984 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3150 9276
rect 3206 9274 3230 9276
rect 3286 9274 3292 9276
rect 3046 9222 3048 9274
rect 3228 9222 3230 9274
rect 2984 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3150 9222
rect 3206 9220 3230 9222
rect 3286 9220 3292 9222
rect 2984 9211 3292 9220
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2288 7644 2596 7653
rect 2288 7642 2294 7644
rect 2350 7642 2374 7644
rect 2430 7642 2454 7644
rect 2510 7642 2534 7644
rect 2590 7642 2596 7644
rect 2350 7590 2352 7642
rect 2532 7590 2534 7642
rect 2288 7588 2294 7590
rect 2350 7588 2374 7590
rect 2430 7588 2454 7590
rect 2510 7588 2534 7590
rect 2590 7588 2596 7590
rect 2288 7579 2596 7588
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 1628 7100 1936 7109
rect 1628 7098 1634 7100
rect 1690 7098 1714 7100
rect 1770 7098 1794 7100
rect 1850 7098 1874 7100
rect 1930 7098 1936 7100
rect 1690 7046 1692 7098
rect 1872 7046 1874 7098
rect 1628 7044 1634 7046
rect 1690 7044 1714 7046
rect 1770 7044 1794 7046
rect 1850 7044 1874 7046
rect 1930 7044 1936 7046
rect 1398 7032 1454 7041
rect 1628 7035 1936 7044
rect 1398 6967 1454 6976
rect 1412 6322 1440 6967
rect 2240 6798 2268 7142
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2136 6792 2188 6798
rect 2228 6792 2280 6798
rect 2136 6734 2188 6740
rect 2226 6760 2228 6769
rect 2280 6760 2282 6769
rect 1596 6458 1624 6734
rect 2056 6458 2084 6734
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1628 6012 1936 6021
rect 1628 6010 1634 6012
rect 1690 6010 1714 6012
rect 1770 6010 1794 6012
rect 1850 6010 1874 6012
rect 1930 6010 1936 6012
rect 1690 5958 1692 6010
rect 1872 5958 1874 6010
rect 1628 5956 1634 5958
rect 1690 5956 1714 5958
rect 1770 5956 1794 5958
rect 1850 5956 1874 5958
rect 1930 5956 1936 5958
rect 1628 5947 1936 5956
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1952 5568 2004 5574
rect 1398 5536 1454 5545
rect 1952 5510 2004 5516
rect 1398 5471 1454 5480
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 938 3360 994 3369
rect 938 3295 994 3304
rect 952 3058 980 3295
rect 940 3052 992 3058
rect 940 2994 992 3000
rect 1320 2990 1348 5170
rect 1628 4924 1936 4933
rect 1628 4922 1634 4924
rect 1690 4922 1714 4924
rect 1770 4922 1794 4924
rect 1850 4922 1874 4924
rect 1930 4922 1936 4924
rect 1690 4870 1692 4922
rect 1872 4870 1874 4922
rect 1628 4868 1634 4870
rect 1690 4868 1714 4870
rect 1770 4868 1794 4870
rect 1850 4868 1874 4870
rect 1930 4868 1936 4870
rect 1628 4859 1936 4868
rect 1964 4622 1992 5510
rect 2056 5098 2084 6258
rect 2148 5370 2176 6734
rect 2608 6730 2636 7414
rect 2700 6905 2728 7686
rect 2792 7002 2820 7754
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2686 6896 2742 6905
rect 2884 6882 2912 8774
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 2984 8188 3292 8197
rect 2984 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3150 8188
rect 3206 8186 3230 8188
rect 3286 8186 3292 8188
rect 3046 8134 3048 8186
rect 3228 8134 3230 8186
rect 2984 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3150 8134
rect 3206 8132 3230 8134
rect 3286 8132 3292 8134
rect 2984 8123 3292 8132
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3252 7290 3280 8026
rect 3344 7954 3372 8230
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3344 7410 3372 7890
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3252 7262 3372 7290
rect 2984 7100 3292 7109
rect 2984 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3150 7100
rect 3206 7098 3230 7100
rect 3286 7098 3292 7100
rect 3046 7046 3048 7098
rect 3228 7046 3230 7098
rect 2984 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3150 7046
rect 3206 7044 3230 7046
rect 3286 7044 3292 7046
rect 2984 7035 3292 7044
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 2884 6866 3004 6882
rect 2884 6860 3016 6866
rect 2884 6854 2964 6860
rect 2686 6831 2742 6840
rect 2964 6802 3016 6808
rect 2226 6695 2282 6704
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2288 6556 2596 6565
rect 2288 6554 2294 6556
rect 2350 6554 2374 6556
rect 2430 6554 2454 6556
rect 2510 6554 2534 6556
rect 2590 6554 2596 6556
rect 2350 6502 2352 6554
rect 2532 6502 2534 6554
rect 2288 6500 2294 6502
rect 2350 6500 2374 6502
rect 2430 6500 2454 6502
rect 2510 6500 2534 6502
rect 2590 6500 2596 6502
rect 2288 6491 2596 6500
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2608 5794 2636 6122
rect 2608 5766 2728 5794
rect 2288 5468 2596 5477
rect 2288 5466 2294 5468
rect 2350 5466 2374 5468
rect 2430 5466 2454 5468
rect 2510 5466 2534 5468
rect 2590 5466 2596 5468
rect 2350 5414 2352 5466
rect 2532 5414 2534 5466
rect 2288 5412 2294 5414
rect 2350 5412 2374 5414
rect 2430 5412 2454 5414
rect 2510 5412 2534 5414
rect 2590 5412 2596 5414
rect 2288 5403 2596 5412
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 4078 1900 4422
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1504 3738 1532 4014
rect 1628 3836 1936 3845
rect 1628 3834 1634 3836
rect 1690 3834 1714 3836
rect 1770 3834 1794 3836
rect 1850 3834 1874 3836
rect 1930 3834 1936 3836
rect 1690 3782 1692 3834
rect 1872 3782 1874 3834
rect 1628 3780 1634 3782
rect 1690 3780 1714 3782
rect 1770 3780 1794 3782
rect 1850 3780 1874 3782
rect 1930 3780 1936 3782
rect 1628 3771 1936 3780
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 3058 1624 3334
rect 2148 3058 2176 5102
rect 2516 4758 2544 5238
rect 2596 5160 2648 5166
rect 2700 5148 2728 5766
rect 2648 5120 2728 5148
rect 2596 5102 2648 5108
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2608 4570 2636 5102
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2700 4729 2728 4966
rect 2686 4720 2742 4729
rect 2686 4655 2742 4664
rect 2608 4542 2728 4570
rect 2288 4380 2596 4389
rect 2288 4378 2294 4380
rect 2350 4378 2374 4380
rect 2430 4378 2454 4380
rect 2510 4378 2534 4380
rect 2590 4378 2596 4380
rect 2350 4326 2352 4378
rect 2532 4326 2534 4378
rect 2288 4324 2294 4326
rect 2350 4324 2374 4326
rect 2430 4324 2454 4326
rect 2510 4324 2534 4326
rect 2590 4324 2596 4326
rect 2288 4315 2596 4324
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2516 3466 2544 4014
rect 2700 3641 2728 4542
rect 2686 3632 2742 3641
rect 2686 3567 2742 3576
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2288 3292 2596 3301
rect 2288 3290 2294 3292
rect 2350 3290 2374 3292
rect 2430 3290 2454 3292
rect 2510 3290 2534 3292
rect 2590 3290 2596 3292
rect 2350 3238 2352 3290
rect 2532 3238 2534 3290
rect 2288 3236 2294 3238
rect 2350 3236 2374 3238
rect 2430 3236 2454 3238
rect 2510 3236 2534 3238
rect 2590 3236 2596 3238
rect 2288 3227 2596 3236
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 2700 2854 2728 3567
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 1628 2748 1936 2757
rect 1628 2746 1634 2748
rect 1690 2746 1714 2748
rect 1770 2746 1794 2748
rect 1850 2746 1874 2748
rect 1930 2746 1936 2748
rect 1690 2694 1692 2746
rect 1872 2694 1874 2746
rect 1628 2692 1634 2694
rect 1690 2692 1714 2694
rect 1770 2692 1794 2694
rect 1850 2692 1874 2694
rect 1930 2692 1936 2694
rect 1628 2683 1936 2692
rect 2288 2204 2596 2213
rect 2288 2202 2294 2204
rect 2350 2202 2374 2204
rect 2430 2202 2454 2204
rect 2510 2202 2534 2204
rect 2590 2202 2596 2204
rect 2350 2150 2352 2202
rect 2532 2150 2534 2202
rect 2288 2148 2294 2150
rect 2350 2148 2374 2150
rect 2430 2148 2454 2150
rect 2510 2148 2534 2150
rect 2590 2148 2596 2150
rect 2288 2139 2596 2148
rect 2792 1465 2820 6258
rect 2884 5302 2912 6598
rect 3160 6118 3188 6938
rect 3240 6792 3292 6798
rect 3344 6780 3372 7262
rect 3436 6798 3464 9318
rect 4264 9110 4292 9590
rect 5368 9574 5488 9602
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 5368 9518 5396 9574
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 4340 9276 4648 9285
rect 4340 9274 4346 9276
rect 4402 9274 4426 9276
rect 4482 9274 4506 9276
rect 4562 9274 4586 9276
rect 4642 9274 4648 9276
rect 4402 9222 4404 9274
rect 4584 9222 4586 9274
rect 4340 9220 4346 9222
rect 4402 9220 4426 9222
rect 4482 9220 4506 9222
rect 4562 9220 4586 9222
rect 4642 9220 4648 9222
rect 4340 9211 4648 9220
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3528 8090 3556 8910
rect 3644 8732 3952 8741
rect 3644 8730 3650 8732
rect 3706 8730 3730 8732
rect 3786 8730 3810 8732
rect 3866 8730 3890 8732
rect 3946 8730 3952 8732
rect 3706 8678 3708 8730
rect 3888 8678 3890 8730
rect 3644 8676 3650 8678
rect 3706 8676 3730 8678
rect 3786 8676 3810 8678
rect 3866 8676 3890 8678
rect 3946 8676 3952 8678
rect 3644 8667 3952 8676
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3644 7644 3952 7653
rect 3644 7642 3650 7644
rect 3706 7642 3730 7644
rect 3786 7642 3810 7644
rect 3866 7642 3890 7644
rect 3946 7642 3952 7644
rect 3706 7590 3708 7642
rect 3888 7590 3890 7642
rect 3644 7588 3650 7590
rect 3706 7588 3730 7590
rect 3786 7588 3810 7590
rect 3866 7588 3890 7590
rect 3946 7588 3952 7590
rect 3644 7579 3952 7588
rect 4080 7546 4108 8910
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3292 6752 3372 6780
rect 3424 6792 3476 6798
rect 3240 6734 3292 6740
rect 3424 6734 3476 6740
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6322 3464 6598
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2984 6012 3292 6021
rect 2984 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3150 6012
rect 3206 6010 3230 6012
rect 3286 6010 3292 6012
rect 3046 5958 3048 6010
rect 3228 5958 3230 6010
rect 2984 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3150 5958
rect 3206 5956 3230 5958
rect 3286 5956 3292 5958
rect 2984 5947 3292 5956
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 3436 5234 3464 6122
rect 3528 5914 3556 7210
rect 3620 7002 3648 7210
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3896 6866 3924 7482
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 4080 6662 4108 7346
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3644 6556 3952 6565
rect 3644 6554 3650 6556
rect 3706 6554 3730 6556
rect 3786 6554 3810 6556
rect 3866 6554 3890 6556
rect 3946 6554 3952 6556
rect 3706 6502 3708 6554
rect 3888 6502 3890 6554
rect 3644 6500 3650 6502
rect 3706 6500 3730 6502
rect 3786 6500 3810 6502
rect 3866 6500 3890 6502
rect 3946 6500 3952 6502
rect 3644 6491 3952 6500
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 4080 5846 4108 6394
rect 4172 6118 4200 8434
rect 4264 7562 4292 8774
rect 4340 8188 4648 8197
rect 4340 8186 4346 8188
rect 4402 8186 4426 8188
rect 4482 8186 4506 8188
rect 4562 8186 4586 8188
rect 4642 8186 4648 8188
rect 4402 8134 4404 8186
rect 4584 8134 4586 8186
rect 4340 8132 4346 8134
rect 4402 8132 4426 8134
rect 4482 8132 4506 8134
rect 4562 8132 4586 8134
rect 4642 8132 4648 8134
rect 4340 8123 4648 8132
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4264 7534 4384 7562
rect 4448 7546 4476 7754
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4264 7002 4292 7414
rect 4356 7206 4384 7534
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4340 7100 4648 7109
rect 4340 7098 4346 7100
rect 4402 7098 4426 7100
rect 4482 7098 4506 7100
rect 4562 7098 4586 7100
rect 4642 7098 4648 7100
rect 4402 7046 4404 7098
rect 4584 7046 4586 7098
rect 4340 7044 4346 7046
rect 4402 7044 4426 7046
rect 4482 7044 4506 7046
rect 4562 7044 4586 7046
rect 4642 7044 4648 7046
rect 4340 7035 4648 7044
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4250 6896 4306 6905
rect 4724 6882 4752 8978
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 8430 4844 8774
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4908 7546 4936 9454
rect 5368 8906 5396 9454
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 9178 5488 9318
rect 5696 9276 6004 9285
rect 5696 9274 5702 9276
rect 5758 9274 5782 9276
rect 5838 9274 5862 9276
rect 5918 9274 5942 9276
rect 5998 9274 6004 9276
rect 5758 9222 5760 9274
rect 5940 9222 5942 9274
rect 5696 9220 5702 9222
rect 5758 9220 5782 9222
rect 5838 9220 5862 9222
rect 5918 9220 5942 9222
rect 5998 9220 6004 9222
rect 5696 9211 6004 9220
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5000 8732 5308 8741
rect 5000 8730 5006 8732
rect 5062 8730 5086 8732
rect 5142 8730 5166 8732
rect 5222 8730 5246 8732
rect 5302 8730 5308 8732
rect 5062 8678 5064 8730
rect 5244 8678 5246 8730
rect 5000 8676 5006 8678
rect 5062 8676 5086 8678
rect 5142 8676 5166 8678
rect 5222 8676 5246 8678
rect 5302 8676 5308 8678
rect 5000 8667 5308 8676
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5000 7818 5028 8502
rect 4988 7812 5040 7818
rect 5040 7772 5396 7800
rect 4988 7754 5040 7760
rect 5000 7644 5308 7653
rect 5000 7642 5006 7644
rect 5062 7642 5086 7644
rect 5142 7642 5166 7644
rect 5222 7642 5246 7644
rect 5302 7642 5308 7644
rect 5062 7590 5064 7642
rect 5244 7590 5246 7642
rect 5000 7588 5006 7590
rect 5062 7588 5086 7590
rect 5142 7588 5166 7590
rect 5222 7588 5246 7590
rect 5302 7588 5308 7590
rect 5000 7579 5308 7588
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4250 6831 4252 6840
rect 4304 6831 4306 6840
rect 4540 6854 4752 6882
rect 4252 6802 4304 6808
rect 4540 6798 4568 6854
rect 4528 6792 4580 6798
rect 4712 6792 4764 6798
rect 4528 6734 4580 6740
rect 4710 6760 4712 6769
rect 4764 6760 4766 6769
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3528 5370 3556 5646
rect 3644 5468 3952 5477
rect 3644 5466 3650 5468
rect 3706 5466 3730 5468
rect 3786 5466 3810 5468
rect 3866 5466 3890 5468
rect 3946 5466 3952 5468
rect 3706 5414 3708 5466
rect 3888 5414 3890 5466
rect 3644 5412 3650 5414
rect 3706 5412 3730 5414
rect 3786 5412 3810 5414
rect 3866 5412 3890 5414
rect 3946 5412 3952 5414
rect 3644 5403 3952 5412
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3528 5234 3556 5306
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 2984 4924 3292 4933
rect 2984 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3150 4924
rect 3206 4922 3230 4924
rect 3286 4922 3292 4924
rect 3046 4870 3048 4922
rect 3228 4870 3230 4922
rect 2984 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3150 4870
rect 3206 4868 3230 4870
rect 3286 4868 3292 4870
rect 2984 4859 3292 4868
rect 2962 4720 3018 4729
rect 2962 4655 3018 4664
rect 2976 4622 3004 4655
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3240 4616 3292 4622
rect 3344 4604 3372 5170
rect 3436 5114 3464 5170
rect 3436 5086 3556 5114
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3292 4576 3372 4604
rect 3240 4558 3292 4564
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 3194 2912 4422
rect 3160 4214 3188 4558
rect 3148 4208 3200 4214
rect 2962 4176 3018 4185
rect 3148 4150 3200 4156
rect 2962 4111 3018 4120
rect 2976 4078 3004 4111
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3252 4010 3280 4558
rect 3436 4146 3464 4966
rect 3528 4690 3556 5086
rect 3988 4826 4016 5646
rect 4080 5302 4108 5782
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4080 4690 4108 5034
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3644 4380 3952 4389
rect 3644 4378 3650 4380
rect 3706 4378 3730 4380
rect 3786 4378 3810 4380
rect 3866 4378 3890 4380
rect 3946 4378 3952 4380
rect 3706 4326 3708 4378
rect 3888 4326 3890 4378
rect 3644 4324 3650 4326
rect 3706 4324 3730 4326
rect 3786 4324 3810 4326
rect 3866 4324 3890 4326
rect 3946 4324 3952 4326
rect 3644 4315 3952 4324
rect 4080 4282 4108 4626
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 2984 3836 3292 3845
rect 2984 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3150 3836
rect 3206 3834 3230 3836
rect 3286 3834 3292 3836
rect 3046 3782 3048 3834
rect 3228 3782 3230 3834
rect 2984 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3150 3782
rect 3206 3780 3230 3782
rect 3286 3780 3292 3782
rect 2984 3771 3292 3780
rect 3344 3466 3372 3878
rect 3528 3720 3556 4218
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3436 3692 3556 3720
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3252 3058 3280 3334
rect 3436 3058 3464 3692
rect 3712 3618 3740 4082
rect 3896 3738 3924 4082
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3528 3590 3740 3618
rect 3528 3194 3556 3590
rect 3644 3292 3952 3301
rect 3644 3290 3650 3292
rect 3706 3290 3730 3292
rect 3786 3290 3810 3292
rect 3866 3290 3890 3292
rect 3946 3290 3952 3292
rect 3706 3238 3708 3290
rect 3888 3238 3890 3290
rect 3644 3236 3650 3238
rect 3706 3236 3730 3238
rect 3786 3236 3810 3238
rect 3866 3236 3890 3238
rect 3946 3236 3952 3238
rect 3644 3227 3952 3236
rect 3988 3194 4016 3946
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 2984 2748 3292 2757
rect 2984 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3150 2748
rect 3206 2746 3230 2748
rect 3286 2746 3292 2748
rect 3046 2694 3048 2746
rect 3228 2694 3230 2746
rect 2984 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3150 2694
rect 3206 2692 3230 2694
rect 3286 2692 3292 2694
rect 2984 2683 3292 2692
rect 3344 2446 3372 2926
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 4080 2378 4108 3878
rect 4172 3534 4200 6054
rect 4264 5846 4292 6666
rect 4540 6254 4568 6734
rect 4710 6695 4766 6704
rect 4724 6390 4752 6695
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4340 6012 4648 6021
rect 4340 6010 4346 6012
rect 4402 6010 4426 6012
rect 4482 6010 4506 6012
rect 4562 6010 4586 6012
rect 4642 6010 4648 6012
rect 4402 5958 4404 6010
rect 4584 5958 4586 6010
rect 4340 5956 4346 5958
rect 4402 5956 4426 5958
rect 4482 5956 4506 5958
rect 4562 5956 4586 5958
rect 4642 5956 4648 5958
rect 4340 5947 4648 5956
rect 4724 5846 4752 6122
rect 4816 5914 4844 7142
rect 4908 6866 4936 7346
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 5092 6798 5120 7278
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 4908 6458 4936 6666
rect 5000 6556 5308 6565
rect 5000 6554 5006 6556
rect 5062 6554 5086 6556
rect 5142 6554 5166 6556
rect 5222 6554 5246 6556
rect 5302 6554 5308 6556
rect 5062 6502 5064 6554
rect 5244 6502 5246 6554
rect 5000 6500 5006 6502
rect 5062 6500 5086 6502
rect 5142 6500 5166 6502
rect 5222 6500 5246 6502
rect 5302 6500 5308 6502
rect 5000 6491 5308 6500
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 5000 5914 5028 6326
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4264 5166 4292 5782
rect 4804 5772 4856 5778
rect 4856 5732 4936 5760
rect 4804 5714 4856 5720
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5370 4752 5510
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4252 5160 4304 5166
rect 4632 5148 4660 5306
rect 4908 5250 4936 5732
rect 5000 5468 5308 5477
rect 5000 5466 5006 5468
rect 5062 5466 5086 5468
rect 5142 5466 5166 5468
rect 5222 5466 5246 5468
rect 5302 5466 5308 5468
rect 5062 5414 5064 5466
rect 5244 5414 5246 5466
rect 5000 5412 5006 5414
rect 5062 5412 5086 5414
rect 5142 5412 5166 5414
rect 5222 5412 5246 5414
rect 5302 5412 5308 5414
rect 5000 5403 5308 5412
rect 5368 5352 5396 7772
rect 5460 7002 5488 9114
rect 6104 9110 6132 9590
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6184 9444 6236 9450
rect 6184 9386 6236 9392
rect 6196 9110 6224 9386
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5696 8188 6004 8197
rect 5696 8186 5702 8188
rect 5758 8186 5782 8188
rect 5838 8186 5862 8188
rect 5918 8186 5942 8188
rect 5998 8186 6004 8188
rect 5758 8134 5760 8186
rect 5940 8134 5942 8186
rect 5696 8132 5702 8134
rect 5758 8132 5782 8134
rect 5838 8132 5862 8134
rect 5918 8132 5942 8134
rect 5998 8132 6004 8134
rect 5696 8123 6004 8132
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5644 7410 5672 8026
rect 6104 7546 6132 8910
rect 6288 8090 6316 9522
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 8809 6776 9318
rect 6734 8800 6790 8809
rect 6356 8732 6664 8741
rect 6734 8735 6790 8744
rect 6356 8730 6362 8732
rect 6418 8730 6442 8732
rect 6498 8730 6522 8732
rect 6578 8730 6602 8732
rect 6658 8730 6664 8732
rect 6418 8678 6420 8730
rect 6600 8678 6602 8730
rect 6356 8676 6362 8678
rect 6418 8676 6442 8678
rect 6498 8676 6522 8678
rect 6578 8676 6602 8678
rect 6658 8676 6664 8678
rect 6356 8667 6664 8676
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6356 7644 6664 7653
rect 6356 7642 6362 7644
rect 6418 7642 6442 7644
rect 6498 7642 6522 7644
rect 6578 7642 6602 7644
rect 6658 7642 6664 7644
rect 6418 7590 6420 7642
rect 6600 7590 6602 7642
rect 6356 7588 6362 7590
rect 6418 7588 6442 7590
rect 6498 7588 6522 7590
rect 6578 7588 6602 7590
rect 6658 7588 6664 7590
rect 6356 7579 6664 7588
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6182 7440 6238 7449
rect 5632 7404 5684 7410
rect 6182 7375 6238 7384
rect 5632 7346 5684 7352
rect 5696 7100 6004 7109
rect 5696 7098 5702 7100
rect 5758 7098 5782 7100
rect 5838 7098 5862 7100
rect 5918 7098 5942 7100
rect 5998 7098 6004 7100
rect 5758 7046 5760 7098
rect 5940 7046 5942 7098
rect 5696 7044 5702 7046
rect 5758 7044 5782 7046
rect 5838 7044 5862 7046
rect 5918 7044 5942 7046
rect 5998 7044 6004 7046
rect 5696 7035 6004 7044
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 6196 6866 6224 7375
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6356 6556 6664 6565
rect 6356 6554 6362 6556
rect 6418 6554 6442 6556
rect 6498 6554 6522 6556
rect 6578 6554 6602 6556
rect 6658 6554 6664 6556
rect 6418 6502 6420 6554
rect 6600 6502 6602 6554
rect 6356 6500 6362 6502
rect 6418 6500 6442 6502
rect 6498 6500 6522 6502
rect 6578 6500 6602 6502
rect 6658 6500 6664 6502
rect 6356 6491 6664 6500
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5276 5324 5396 5352
rect 4908 5234 5028 5250
rect 4908 5228 5040 5234
rect 4908 5222 4988 5228
rect 4988 5170 5040 5176
rect 4632 5120 4752 5148
rect 4252 5102 4304 5108
rect 4340 4924 4648 4933
rect 4340 4922 4346 4924
rect 4402 4922 4426 4924
rect 4482 4922 4506 4924
rect 4562 4922 4586 4924
rect 4642 4922 4648 4924
rect 4402 4870 4404 4922
rect 4584 4870 4586 4922
rect 4340 4868 4346 4870
rect 4402 4868 4426 4870
rect 4482 4868 4506 4870
rect 4562 4868 4586 4870
rect 4642 4868 4648 4870
rect 4340 4859 4648 4868
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4264 3058 4292 4422
rect 4356 4078 4384 4558
rect 4724 4214 4752 5120
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4340 3836 4648 3845
rect 4340 3834 4346 3836
rect 4402 3834 4426 3836
rect 4482 3834 4506 3836
rect 4562 3834 4586 3836
rect 4642 3834 4648 3836
rect 4402 3782 4404 3834
rect 4584 3782 4586 3834
rect 4340 3780 4346 3782
rect 4402 3780 4426 3782
rect 4482 3780 4506 3782
rect 4562 3780 4586 3782
rect 4642 3780 4648 3782
rect 4340 3771 4648 3780
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4540 3058 4568 3674
rect 4724 3194 4752 4014
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4816 2922 4844 5034
rect 5000 4690 5028 5034
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5276 4554 5304 5324
rect 5460 5166 5488 6394
rect 6092 6112 6144 6118
rect 6090 6080 6092 6089
rect 6144 6080 6146 6089
rect 5696 6012 6004 6021
rect 6090 6015 6146 6024
rect 5696 6010 5702 6012
rect 5758 6010 5782 6012
rect 5838 6010 5862 6012
rect 5918 6010 5942 6012
rect 5998 6010 6004 6012
rect 5758 5958 5760 6010
rect 5940 5958 5942 6010
rect 5696 5956 5702 5958
rect 5758 5956 5782 5958
rect 5838 5956 5862 5958
rect 5918 5956 5942 5958
rect 5998 5956 6004 5958
rect 5696 5947 6004 5956
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5264 4548 5316 4554
rect 4908 4508 5264 4536
rect 4908 4214 4936 4508
rect 5264 4490 5316 4496
rect 5000 4380 5308 4389
rect 5000 4378 5006 4380
rect 5062 4378 5086 4380
rect 5142 4378 5166 4380
rect 5222 4378 5246 4380
rect 5302 4378 5308 4380
rect 5062 4326 5064 4378
rect 5244 4326 5246 4378
rect 5000 4324 5006 4326
rect 5062 4324 5086 4326
rect 5142 4324 5166 4326
rect 5222 4324 5246 4326
rect 5302 4324 5308 4326
rect 5000 4315 5308 4324
rect 4896 4208 4948 4214
rect 4894 4176 4896 4185
rect 4948 4176 4950 4185
rect 4894 4111 4950 4120
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5092 3738 5120 3878
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5000 3292 5308 3301
rect 5000 3290 5006 3292
rect 5062 3290 5086 3292
rect 5142 3290 5166 3292
rect 5222 3290 5246 3292
rect 5302 3290 5308 3292
rect 5062 3238 5064 3290
rect 5244 3238 5246 3290
rect 5000 3236 5006 3238
rect 5062 3236 5086 3238
rect 5142 3236 5166 3238
rect 5222 3236 5246 3238
rect 5302 3236 5308 3238
rect 5000 3227 5308 3236
rect 5368 3058 5396 5034
rect 5460 3602 5488 5102
rect 5552 3738 5580 5238
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 5696 4924 6004 4933
rect 5696 4922 5702 4924
rect 5758 4922 5782 4924
rect 5838 4922 5862 4924
rect 5918 4922 5942 4924
rect 5998 4922 6004 4924
rect 5758 4870 5760 4922
rect 5940 4870 5942 4922
rect 5696 4868 5702 4870
rect 5758 4868 5782 4870
rect 5838 4868 5862 4870
rect 5918 4868 5942 4870
rect 5998 4868 6004 4870
rect 5696 4859 6004 4868
rect 6104 3942 6132 5170
rect 6196 4729 6224 5510
rect 6288 4826 6316 5578
rect 6356 5468 6664 5477
rect 6356 5466 6362 5468
rect 6418 5466 6442 5468
rect 6498 5466 6522 5468
rect 6578 5466 6602 5468
rect 6658 5466 6664 5468
rect 6418 5414 6420 5466
rect 6600 5414 6602 5466
rect 6356 5412 6362 5414
rect 6418 5412 6442 5414
rect 6498 5412 6522 5414
rect 6578 5412 6602 5414
rect 6658 5412 6664 5414
rect 6356 5403 6664 5412
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6182 4720 6238 4729
rect 6182 4655 6238 4664
rect 6288 4604 6316 4762
rect 6196 4576 6316 4604
rect 6196 4486 6224 4576
rect 6380 4536 6408 4966
rect 6288 4508 6408 4536
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 5696 3836 6004 3845
rect 5696 3834 5702 3836
rect 5758 3834 5782 3836
rect 5838 3834 5862 3836
rect 5918 3834 5942 3836
rect 5998 3834 6004 3836
rect 5758 3782 5760 3834
rect 5940 3782 5942 3834
rect 5696 3780 5702 3782
rect 5758 3780 5782 3782
rect 5838 3780 5862 3782
rect 5918 3780 5942 3782
rect 5998 3780 6004 3782
rect 5696 3771 6004 3780
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5828 3641 5856 3674
rect 5814 3632 5870 3641
rect 5448 3596 5500 3602
rect 5814 3567 5870 3576
rect 5448 3538 5500 3544
rect 6104 3058 6132 3878
rect 6196 3534 6224 4422
rect 6288 3738 6316 4508
rect 6356 4380 6664 4389
rect 6356 4378 6362 4380
rect 6418 4378 6442 4380
rect 6498 4378 6522 4380
rect 6578 4378 6602 4380
rect 6658 4378 6664 4380
rect 6418 4326 6420 4378
rect 6600 4326 6602 4378
rect 6356 4324 6362 4326
rect 6418 4324 6442 4326
rect 6498 4324 6522 4326
rect 6578 4324 6602 4326
rect 6658 4324 6664 4326
rect 6356 4315 6664 4324
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6734 3360 6790 3369
rect 6356 3292 6664 3301
rect 6734 3295 6790 3304
rect 6356 3290 6362 3292
rect 6418 3290 6442 3292
rect 6498 3290 6522 3292
rect 6578 3290 6602 3292
rect 6658 3290 6664 3292
rect 6418 3238 6420 3290
rect 6600 3238 6602 3290
rect 6356 3236 6362 3238
rect 6418 3236 6442 3238
rect 6498 3236 6522 3238
rect 6578 3236 6602 3238
rect 6658 3236 6664 3238
rect 6356 3227 6664 3236
rect 6748 3194 6776 3295
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 4340 2748 4648 2757
rect 4340 2746 4346 2748
rect 4402 2746 4426 2748
rect 4482 2746 4506 2748
rect 4562 2746 4586 2748
rect 4642 2746 4648 2748
rect 4402 2694 4404 2746
rect 4584 2694 4586 2746
rect 4340 2692 4346 2694
rect 4402 2692 4426 2694
rect 4482 2692 4506 2694
rect 4562 2692 4586 2694
rect 4642 2692 4648 2694
rect 4340 2683 4648 2692
rect 5696 2748 6004 2757
rect 5696 2746 5702 2748
rect 5758 2746 5782 2748
rect 5838 2746 5862 2748
rect 5918 2746 5942 2748
rect 5998 2746 6004 2748
rect 5758 2694 5760 2746
rect 5940 2694 5942 2746
rect 5696 2692 5702 2694
rect 5758 2692 5782 2694
rect 5838 2692 5862 2694
rect 5918 2692 5942 2694
rect 5998 2692 6004 2694
rect 5696 2683 6004 2692
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 3644 2204 3952 2213
rect 3644 2202 3650 2204
rect 3706 2202 3730 2204
rect 3786 2202 3810 2204
rect 3866 2202 3890 2204
rect 3946 2202 3952 2204
rect 3706 2150 3708 2202
rect 3888 2150 3890 2202
rect 3644 2148 3650 2150
rect 3706 2148 3730 2150
rect 3786 2148 3810 2150
rect 3866 2148 3890 2150
rect 3946 2148 3952 2150
rect 3644 2139 3952 2148
rect 5000 2204 5308 2213
rect 5000 2202 5006 2204
rect 5062 2202 5086 2204
rect 5142 2202 5166 2204
rect 5222 2202 5246 2204
rect 5302 2202 5308 2204
rect 5062 2150 5064 2202
rect 5244 2150 5246 2202
rect 5000 2148 5006 2150
rect 5062 2148 5086 2150
rect 5142 2148 5166 2150
rect 5222 2148 5246 2150
rect 5302 2148 5308 2150
rect 5000 2139 5308 2148
rect 5552 2009 5580 2246
rect 5538 2000 5594 2009
rect 5538 1935 5594 1944
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 6196 649 6224 2246
rect 6356 2204 6664 2213
rect 6356 2202 6362 2204
rect 6418 2202 6442 2204
rect 6498 2202 6522 2204
rect 6578 2202 6602 2204
rect 6658 2202 6664 2204
rect 6418 2150 6420 2202
rect 6600 2150 6602 2202
rect 6356 2148 6362 2150
rect 6418 2148 6442 2150
rect 6498 2148 6522 2150
rect 6578 2148 6602 2150
rect 6658 2148 6664 2150
rect 6356 2139 6664 2148
rect 6182 640 6238 649
rect 6182 575 6238 584
<< via2 >>
rect 6366 11464 6422 11520
rect 938 10920 994 10976
rect 1634 10362 1690 10364
rect 1714 10362 1770 10364
rect 1794 10362 1850 10364
rect 1874 10362 1930 10364
rect 1634 10310 1680 10362
rect 1680 10310 1690 10362
rect 1714 10310 1744 10362
rect 1744 10310 1756 10362
rect 1756 10310 1770 10362
rect 1794 10310 1808 10362
rect 1808 10310 1820 10362
rect 1820 10310 1850 10362
rect 1874 10310 1884 10362
rect 1884 10310 1930 10362
rect 1634 10308 1690 10310
rect 1714 10308 1770 10310
rect 1794 10308 1850 10310
rect 1874 10308 1930 10310
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 3150 10362 3206 10364
rect 3230 10362 3286 10364
rect 2990 10310 3036 10362
rect 3036 10310 3046 10362
rect 3070 10310 3100 10362
rect 3100 10310 3112 10362
rect 3112 10310 3126 10362
rect 3150 10310 3164 10362
rect 3164 10310 3176 10362
rect 3176 10310 3206 10362
rect 3230 10310 3240 10362
rect 3240 10310 3286 10362
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 3150 10308 3206 10310
rect 3230 10308 3286 10310
rect 4346 10362 4402 10364
rect 4426 10362 4482 10364
rect 4506 10362 4562 10364
rect 4586 10362 4642 10364
rect 4346 10310 4392 10362
rect 4392 10310 4402 10362
rect 4426 10310 4456 10362
rect 4456 10310 4468 10362
rect 4468 10310 4482 10362
rect 4506 10310 4520 10362
rect 4520 10310 4532 10362
rect 4532 10310 4562 10362
rect 4586 10310 4596 10362
rect 4596 10310 4642 10362
rect 4346 10308 4402 10310
rect 4426 10308 4482 10310
rect 4506 10308 4562 10310
rect 4586 10308 4642 10310
rect 5702 10362 5758 10364
rect 5782 10362 5838 10364
rect 5862 10362 5918 10364
rect 5942 10362 5998 10364
rect 5702 10310 5748 10362
rect 5748 10310 5758 10362
rect 5782 10310 5812 10362
rect 5812 10310 5824 10362
rect 5824 10310 5838 10362
rect 5862 10310 5876 10362
rect 5876 10310 5888 10362
rect 5888 10310 5918 10362
rect 5942 10310 5952 10362
rect 5952 10310 5998 10362
rect 5702 10308 5758 10310
rect 5782 10308 5838 10310
rect 5862 10308 5918 10310
rect 5942 10308 5998 10310
rect 5354 10104 5410 10160
rect 2294 9818 2350 9820
rect 2374 9818 2430 9820
rect 2454 9818 2510 9820
rect 2534 9818 2590 9820
rect 2294 9766 2340 9818
rect 2340 9766 2350 9818
rect 2374 9766 2404 9818
rect 2404 9766 2416 9818
rect 2416 9766 2430 9818
rect 2454 9766 2468 9818
rect 2468 9766 2480 9818
rect 2480 9766 2510 9818
rect 2534 9766 2544 9818
rect 2544 9766 2590 9818
rect 2294 9764 2350 9766
rect 2374 9764 2430 9766
rect 2454 9764 2510 9766
rect 2534 9764 2590 9766
rect 1634 9274 1690 9276
rect 1714 9274 1770 9276
rect 1794 9274 1850 9276
rect 1874 9274 1930 9276
rect 1634 9222 1680 9274
rect 1680 9222 1690 9274
rect 1714 9222 1744 9274
rect 1744 9222 1756 9274
rect 1756 9222 1770 9274
rect 1794 9222 1808 9274
rect 1808 9222 1820 9274
rect 1820 9222 1850 9274
rect 1874 9222 1884 9274
rect 1884 9222 1930 9274
rect 1634 9220 1690 9222
rect 1714 9220 1770 9222
rect 1794 9220 1850 9222
rect 1874 9220 1930 9222
rect 938 9016 994 9072
rect 2294 8730 2350 8732
rect 2374 8730 2430 8732
rect 2454 8730 2510 8732
rect 2534 8730 2590 8732
rect 2294 8678 2340 8730
rect 2340 8678 2350 8730
rect 2374 8678 2404 8730
rect 2404 8678 2416 8730
rect 2416 8678 2430 8730
rect 2454 8678 2468 8730
rect 2468 8678 2480 8730
rect 2480 8678 2510 8730
rect 2534 8678 2544 8730
rect 2544 8678 2590 8730
rect 2294 8676 2350 8678
rect 2374 8676 2430 8678
rect 2454 8676 2510 8678
rect 2534 8676 2590 8678
rect 1634 8186 1690 8188
rect 1714 8186 1770 8188
rect 1794 8186 1850 8188
rect 1874 8186 1930 8188
rect 1634 8134 1680 8186
rect 1680 8134 1690 8186
rect 1714 8134 1744 8186
rect 1744 8134 1756 8186
rect 1756 8134 1770 8186
rect 1794 8134 1808 8186
rect 1808 8134 1820 8186
rect 1820 8134 1850 8186
rect 1874 8134 1884 8186
rect 1884 8134 1930 8186
rect 1634 8132 1690 8134
rect 1714 8132 1770 8134
rect 1794 8132 1850 8134
rect 1874 8132 1930 8134
rect 3650 9818 3706 9820
rect 3730 9818 3786 9820
rect 3810 9818 3866 9820
rect 3890 9818 3946 9820
rect 3650 9766 3696 9818
rect 3696 9766 3706 9818
rect 3730 9766 3760 9818
rect 3760 9766 3772 9818
rect 3772 9766 3786 9818
rect 3810 9766 3824 9818
rect 3824 9766 3836 9818
rect 3836 9766 3866 9818
rect 3890 9766 3900 9818
rect 3900 9766 3946 9818
rect 3650 9764 3706 9766
rect 3730 9764 3786 9766
rect 3810 9764 3866 9766
rect 3890 9764 3946 9766
rect 5006 9818 5062 9820
rect 5086 9818 5142 9820
rect 5166 9818 5222 9820
rect 5246 9818 5302 9820
rect 5006 9766 5052 9818
rect 5052 9766 5062 9818
rect 5086 9766 5116 9818
rect 5116 9766 5128 9818
rect 5128 9766 5142 9818
rect 5166 9766 5180 9818
rect 5180 9766 5192 9818
rect 5192 9766 5222 9818
rect 5246 9766 5256 9818
rect 5256 9766 5302 9818
rect 5006 9764 5062 9766
rect 5086 9764 5142 9766
rect 5166 9764 5222 9766
rect 5246 9764 5302 9766
rect 6362 9818 6418 9820
rect 6442 9818 6498 9820
rect 6522 9818 6578 9820
rect 6602 9818 6658 9820
rect 6362 9766 6408 9818
rect 6408 9766 6418 9818
rect 6442 9766 6472 9818
rect 6472 9766 6484 9818
rect 6484 9766 6498 9818
rect 6522 9766 6536 9818
rect 6536 9766 6548 9818
rect 6548 9766 6578 9818
rect 6602 9766 6612 9818
rect 6612 9766 6658 9818
rect 6362 9764 6418 9766
rect 6442 9764 6498 9766
rect 6522 9764 6578 9766
rect 6602 9764 6658 9766
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 3150 9274 3206 9276
rect 3230 9274 3286 9276
rect 2990 9222 3036 9274
rect 3036 9222 3046 9274
rect 3070 9222 3100 9274
rect 3100 9222 3112 9274
rect 3112 9222 3126 9274
rect 3150 9222 3164 9274
rect 3164 9222 3176 9274
rect 3176 9222 3206 9274
rect 3230 9222 3240 9274
rect 3240 9222 3286 9274
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 3150 9220 3206 9222
rect 3230 9220 3286 9222
rect 2294 7642 2350 7644
rect 2374 7642 2430 7644
rect 2454 7642 2510 7644
rect 2534 7642 2590 7644
rect 2294 7590 2340 7642
rect 2340 7590 2350 7642
rect 2374 7590 2404 7642
rect 2404 7590 2416 7642
rect 2416 7590 2430 7642
rect 2454 7590 2468 7642
rect 2468 7590 2480 7642
rect 2480 7590 2510 7642
rect 2534 7590 2544 7642
rect 2544 7590 2590 7642
rect 2294 7588 2350 7590
rect 2374 7588 2430 7590
rect 2454 7588 2510 7590
rect 2534 7588 2590 7590
rect 1634 7098 1690 7100
rect 1714 7098 1770 7100
rect 1794 7098 1850 7100
rect 1874 7098 1930 7100
rect 1634 7046 1680 7098
rect 1680 7046 1690 7098
rect 1714 7046 1744 7098
rect 1744 7046 1756 7098
rect 1756 7046 1770 7098
rect 1794 7046 1808 7098
rect 1808 7046 1820 7098
rect 1820 7046 1850 7098
rect 1874 7046 1884 7098
rect 1884 7046 1930 7098
rect 1634 7044 1690 7046
rect 1714 7044 1770 7046
rect 1794 7044 1850 7046
rect 1874 7044 1930 7046
rect 1398 6976 1454 7032
rect 2226 6740 2228 6760
rect 2228 6740 2280 6760
rect 2280 6740 2282 6760
rect 1634 6010 1690 6012
rect 1714 6010 1770 6012
rect 1794 6010 1850 6012
rect 1874 6010 1930 6012
rect 1634 5958 1680 6010
rect 1680 5958 1690 6010
rect 1714 5958 1744 6010
rect 1744 5958 1756 6010
rect 1756 5958 1770 6010
rect 1794 5958 1808 6010
rect 1808 5958 1820 6010
rect 1820 5958 1850 6010
rect 1874 5958 1884 6010
rect 1884 5958 1930 6010
rect 1634 5956 1690 5958
rect 1714 5956 1770 5958
rect 1794 5956 1850 5958
rect 1874 5956 1930 5958
rect 1398 5480 1454 5536
rect 938 3304 994 3360
rect 1634 4922 1690 4924
rect 1714 4922 1770 4924
rect 1794 4922 1850 4924
rect 1874 4922 1930 4924
rect 1634 4870 1680 4922
rect 1680 4870 1690 4922
rect 1714 4870 1744 4922
rect 1744 4870 1756 4922
rect 1756 4870 1770 4922
rect 1794 4870 1808 4922
rect 1808 4870 1820 4922
rect 1820 4870 1850 4922
rect 1874 4870 1884 4922
rect 1884 4870 1930 4922
rect 1634 4868 1690 4870
rect 1714 4868 1770 4870
rect 1794 4868 1850 4870
rect 1874 4868 1930 4870
rect 2226 6704 2282 6740
rect 2686 6840 2742 6896
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 3150 8186 3206 8188
rect 3230 8186 3286 8188
rect 2990 8134 3036 8186
rect 3036 8134 3046 8186
rect 3070 8134 3100 8186
rect 3100 8134 3112 8186
rect 3112 8134 3126 8186
rect 3150 8134 3164 8186
rect 3164 8134 3176 8186
rect 3176 8134 3206 8186
rect 3230 8134 3240 8186
rect 3240 8134 3286 8186
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 3150 8132 3206 8134
rect 3230 8132 3286 8134
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 3150 7098 3206 7100
rect 3230 7098 3286 7100
rect 2990 7046 3036 7098
rect 3036 7046 3046 7098
rect 3070 7046 3100 7098
rect 3100 7046 3112 7098
rect 3112 7046 3126 7098
rect 3150 7046 3164 7098
rect 3164 7046 3176 7098
rect 3176 7046 3206 7098
rect 3230 7046 3240 7098
rect 3240 7046 3286 7098
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 3150 7044 3206 7046
rect 3230 7044 3286 7046
rect 2294 6554 2350 6556
rect 2374 6554 2430 6556
rect 2454 6554 2510 6556
rect 2534 6554 2590 6556
rect 2294 6502 2340 6554
rect 2340 6502 2350 6554
rect 2374 6502 2404 6554
rect 2404 6502 2416 6554
rect 2416 6502 2430 6554
rect 2454 6502 2468 6554
rect 2468 6502 2480 6554
rect 2480 6502 2510 6554
rect 2534 6502 2544 6554
rect 2544 6502 2590 6554
rect 2294 6500 2350 6502
rect 2374 6500 2430 6502
rect 2454 6500 2510 6502
rect 2534 6500 2590 6502
rect 2294 5466 2350 5468
rect 2374 5466 2430 5468
rect 2454 5466 2510 5468
rect 2534 5466 2590 5468
rect 2294 5414 2340 5466
rect 2340 5414 2350 5466
rect 2374 5414 2404 5466
rect 2404 5414 2416 5466
rect 2416 5414 2430 5466
rect 2454 5414 2468 5466
rect 2468 5414 2480 5466
rect 2480 5414 2510 5466
rect 2534 5414 2544 5466
rect 2544 5414 2590 5466
rect 2294 5412 2350 5414
rect 2374 5412 2430 5414
rect 2454 5412 2510 5414
rect 2534 5412 2590 5414
rect 1634 3834 1690 3836
rect 1714 3834 1770 3836
rect 1794 3834 1850 3836
rect 1874 3834 1930 3836
rect 1634 3782 1680 3834
rect 1680 3782 1690 3834
rect 1714 3782 1744 3834
rect 1744 3782 1756 3834
rect 1756 3782 1770 3834
rect 1794 3782 1808 3834
rect 1808 3782 1820 3834
rect 1820 3782 1850 3834
rect 1874 3782 1884 3834
rect 1884 3782 1930 3834
rect 1634 3780 1690 3782
rect 1714 3780 1770 3782
rect 1794 3780 1850 3782
rect 1874 3780 1930 3782
rect 2686 4664 2742 4720
rect 2294 4378 2350 4380
rect 2374 4378 2430 4380
rect 2454 4378 2510 4380
rect 2534 4378 2590 4380
rect 2294 4326 2340 4378
rect 2340 4326 2350 4378
rect 2374 4326 2404 4378
rect 2404 4326 2416 4378
rect 2416 4326 2430 4378
rect 2454 4326 2468 4378
rect 2468 4326 2480 4378
rect 2480 4326 2510 4378
rect 2534 4326 2544 4378
rect 2544 4326 2590 4378
rect 2294 4324 2350 4326
rect 2374 4324 2430 4326
rect 2454 4324 2510 4326
rect 2534 4324 2590 4326
rect 2686 3576 2742 3632
rect 2294 3290 2350 3292
rect 2374 3290 2430 3292
rect 2454 3290 2510 3292
rect 2534 3290 2590 3292
rect 2294 3238 2340 3290
rect 2340 3238 2350 3290
rect 2374 3238 2404 3290
rect 2404 3238 2416 3290
rect 2416 3238 2430 3290
rect 2454 3238 2468 3290
rect 2468 3238 2480 3290
rect 2480 3238 2510 3290
rect 2534 3238 2544 3290
rect 2544 3238 2590 3290
rect 2294 3236 2350 3238
rect 2374 3236 2430 3238
rect 2454 3236 2510 3238
rect 2534 3236 2590 3238
rect 1634 2746 1690 2748
rect 1714 2746 1770 2748
rect 1794 2746 1850 2748
rect 1874 2746 1930 2748
rect 1634 2694 1680 2746
rect 1680 2694 1690 2746
rect 1714 2694 1744 2746
rect 1744 2694 1756 2746
rect 1756 2694 1770 2746
rect 1794 2694 1808 2746
rect 1808 2694 1820 2746
rect 1820 2694 1850 2746
rect 1874 2694 1884 2746
rect 1884 2694 1930 2746
rect 1634 2692 1690 2694
rect 1714 2692 1770 2694
rect 1794 2692 1850 2694
rect 1874 2692 1930 2694
rect 2294 2202 2350 2204
rect 2374 2202 2430 2204
rect 2454 2202 2510 2204
rect 2534 2202 2590 2204
rect 2294 2150 2340 2202
rect 2340 2150 2350 2202
rect 2374 2150 2404 2202
rect 2404 2150 2416 2202
rect 2416 2150 2430 2202
rect 2454 2150 2468 2202
rect 2468 2150 2480 2202
rect 2480 2150 2510 2202
rect 2534 2150 2544 2202
rect 2544 2150 2590 2202
rect 2294 2148 2350 2150
rect 2374 2148 2430 2150
rect 2454 2148 2510 2150
rect 2534 2148 2590 2150
rect 4346 9274 4402 9276
rect 4426 9274 4482 9276
rect 4506 9274 4562 9276
rect 4586 9274 4642 9276
rect 4346 9222 4392 9274
rect 4392 9222 4402 9274
rect 4426 9222 4456 9274
rect 4456 9222 4468 9274
rect 4468 9222 4482 9274
rect 4506 9222 4520 9274
rect 4520 9222 4532 9274
rect 4532 9222 4562 9274
rect 4586 9222 4596 9274
rect 4596 9222 4642 9274
rect 4346 9220 4402 9222
rect 4426 9220 4482 9222
rect 4506 9220 4562 9222
rect 4586 9220 4642 9222
rect 3650 8730 3706 8732
rect 3730 8730 3786 8732
rect 3810 8730 3866 8732
rect 3890 8730 3946 8732
rect 3650 8678 3696 8730
rect 3696 8678 3706 8730
rect 3730 8678 3760 8730
rect 3760 8678 3772 8730
rect 3772 8678 3786 8730
rect 3810 8678 3824 8730
rect 3824 8678 3836 8730
rect 3836 8678 3866 8730
rect 3890 8678 3900 8730
rect 3900 8678 3946 8730
rect 3650 8676 3706 8678
rect 3730 8676 3786 8678
rect 3810 8676 3866 8678
rect 3890 8676 3946 8678
rect 3650 7642 3706 7644
rect 3730 7642 3786 7644
rect 3810 7642 3866 7644
rect 3890 7642 3946 7644
rect 3650 7590 3696 7642
rect 3696 7590 3706 7642
rect 3730 7590 3760 7642
rect 3760 7590 3772 7642
rect 3772 7590 3786 7642
rect 3810 7590 3824 7642
rect 3824 7590 3836 7642
rect 3836 7590 3866 7642
rect 3890 7590 3900 7642
rect 3900 7590 3946 7642
rect 3650 7588 3706 7590
rect 3730 7588 3786 7590
rect 3810 7588 3866 7590
rect 3890 7588 3946 7590
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 3150 6010 3206 6012
rect 3230 6010 3286 6012
rect 2990 5958 3036 6010
rect 3036 5958 3046 6010
rect 3070 5958 3100 6010
rect 3100 5958 3112 6010
rect 3112 5958 3126 6010
rect 3150 5958 3164 6010
rect 3164 5958 3176 6010
rect 3176 5958 3206 6010
rect 3230 5958 3240 6010
rect 3240 5958 3286 6010
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 3150 5956 3206 5958
rect 3230 5956 3286 5958
rect 3650 6554 3706 6556
rect 3730 6554 3786 6556
rect 3810 6554 3866 6556
rect 3890 6554 3946 6556
rect 3650 6502 3696 6554
rect 3696 6502 3706 6554
rect 3730 6502 3760 6554
rect 3760 6502 3772 6554
rect 3772 6502 3786 6554
rect 3810 6502 3824 6554
rect 3824 6502 3836 6554
rect 3836 6502 3866 6554
rect 3890 6502 3900 6554
rect 3900 6502 3946 6554
rect 3650 6500 3706 6502
rect 3730 6500 3786 6502
rect 3810 6500 3866 6502
rect 3890 6500 3946 6502
rect 4346 8186 4402 8188
rect 4426 8186 4482 8188
rect 4506 8186 4562 8188
rect 4586 8186 4642 8188
rect 4346 8134 4392 8186
rect 4392 8134 4402 8186
rect 4426 8134 4456 8186
rect 4456 8134 4468 8186
rect 4468 8134 4482 8186
rect 4506 8134 4520 8186
rect 4520 8134 4532 8186
rect 4532 8134 4562 8186
rect 4586 8134 4596 8186
rect 4596 8134 4642 8186
rect 4346 8132 4402 8134
rect 4426 8132 4482 8134
rect 4506 8132 4562 8134
rect 4586 8132 4642 8134
rect 4346 7098 4402 7100
rect 4426 7098 4482 7100
rect 4506 7098 4562 7100
rect 4586 7098 4642 7100
rect 4346 7046 4392 7098
rect 4392 7046 4402 7098
rect 4426 7046 4456 7098
rect 4456 7046 4468 7098
rect 4468 7046 4482 7098
rect 4506 7046 4520 7098
rect 4520 7046 4532 7098
rect 4532 7046 4562 7098
rect 4586 7046 4596 7098
rect 4596 7046 4642 7098
rect 4346 7044 4402 7046
rect 4426 7044 4482 7046
rect 4506 7044 4562 7046
rect 4586 7044 4642 7046
rect 4250 6860 4306 6896
rect 5702 9274 5758 9276
rect 5782 9274 5838 9276
rect 5862 9274 5918 9276
rect 5942 9274 5998 9276
rect 5702 9222 5748 9274
rect 5748 9222 5758 9274
rect 5782 9222 5812 9274
rect 5812 9222 5824 9274
rect 5824 9222 5838 9274
rect 5862 9222 5876 9274
rect 5876 9222 5888 9274
rect 5888 9222 5918 9274
rect 5942 9222 5952 9274
rect 5952 9222 5998 9274
rect 5702 9220 5758 9222
rect 5782 9220 5838 9222
rect 5862 9220 5918 9222
rect 5942 9220 5998 9222
rect 5006 8730 5062 8732
rect 5086 8730 5142 8732
rect 5166 8730 5222 8732
rect 5246 8730 5302 8732
rect 5006 8678 5052 8730
rect 5052 8678 5062 8730
rect 5086 8678 5116 8730
rect 5116 8678 5128 8730
rect 5128 8678 5142 8730
rect 5166 8678 5180 8730
rect 5180 8678 5192 8730
rect 5192 8678 5222 8730
rect 5246 8678 5256 8730
rect 5256 8678 5302 8730
rect 5006 8676 5062 8678
rect 5086 8676 5142 8678
rect 5166 8676 5222 8678
rect 5246 8676 5302 8678
rect 5006 7642 5062 7644
rect 5086 7642 5142 7644
rect 5166 7642 5222 7644
rect 5246 7642 5302 7644
rect 5006 7590 5052 7642
rect 5052 7590 5062 7642
rect 5086 7590 5116 7642
rect 5116 7590 5128 7642
rect 5128 7590 5142 7642
rect 5166 7590 5180 7642
rect 5180 7590 5192 7642
rect 5192 7590 5222 7642
rect 5246 7590 5256 7642
rect 5256 7590 5302 7642
rect 5006 7588 5062 7590
rect 5086 7588 5142 7590
rect 5166 7588 5222 7590
rect 5246 7588 5302 7590
rect 4250 6840 4252 6860
rect 4252 6840 4304 6860
rect 4304 6840 4306 6860
rect 4710 6740 4712 6760
rect 4712 6740 4764 6760
rect 4764 6740 4766 6760
rect 3650 5466 3706 5468
rect 3730 5466 3786 5468
rect 3810 5466 3866 5468
rect 3890 5466 3946 5468
rect 3650 5414 3696 5466
rect 3696 5414 3706 5466
rect 3730 5414 3760 5466
rect 3760 5414 3772 5466
rect 3772 5414 3786 5466
rect 3810 5414 3824 5466
rect 3824 5414 3836 5466
rect 3836 5414 3866 5466
rect 3890 5414 3900 5466
rect 3900 5414 3946 5466
rect 3650 5412 3706 5414
rect 3730 5412 3786 5414
rect 3810 5412 3866 5414
rect 3890 5412 3946 5414
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 3150 4922 3206 4924
rect 3230 4922 3286 4924
rect 2990 4870 3036 4922
rect 3036 4870 3046 4922
rect 3070 4870 3100 4922
rect 3100 4870 3112 4922
rect 3112 4870 3126 4922
rect 3150 4870 3164 4922
rect 3164 4870 3176 4922
rect 3176 4870 3206 4922
rect 3230 4870 3240 4922
rect 3240 4870 3286 4922
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 3150 4868 3206 4870
rect 3230 4868 3286 4870
rect 2962 4664 3018 4720
rect 2962 4120 3018 4176
rect 3650 4378 3706 4380
rect 3730 4378 3786 4380
rect 3810 4378 3866 4380
rect 3890 4378 3946 4380
rect 3650 4326 3696 4378
rect 3696 4326 3706 4378
rect 3730 4326 3760 4378
rect 3760 4326 3772 4378
rect 3772 4326 3786 4378
rect 3810 4326 3824 4378
rect 3824 4326 3836 4378
rect 3836 4326 3866 4378
rect 3890 4326 3900 4378
rect 3900 4326 3946 4378
rect 3650 4324 3706 4326
rect 3730 4324 3786 4326
rect 3810 4324 3866 4326
rect 3890 4324 3946 4326
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 3150 3834 3206 3836
rect 3230 3834 3286 3836
rect 2990 3782 3036 3834
rect 3036 3782 3046 3834
rect 3070 3782 3100 3834
rect 3100 3782 3112 3834
rect 3112 3782 3126 3834
rect 3150 3782 3164 3834
rect 3164 3782 3176 3834
rect 3176 3782 3206 3834
rect 3230 3782 3240 3834
rect 3240 3782 3286 3834
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 3150 3780 3206 3782
rect 3230 3780 3286 3782
rect 3650 3290 3706 3292
rect 3730 3290 3786 3292
rect 3810 3290 3866 3292
rect 3890 3290 3946 3292
rect 3650 3238 3696 3290
rect 3696 3238 3706 3290
rect 3730 3238 3760 3290
rect 3760 3238 3772 3290
rect 3772 3238 3786 3290
rect 3810 3238 3824 3290
rect 3824 3238 3836 3290
rect 3836 3238 3866 3290
rect 3890 3238 3900 3290
rect 3900 3238 3946 3290
rect 3650 3236 3706 3238
rect 3730 3236 3786 3238
rect 3810 3236 3866 3238
rect 3890 3236 3946 3238
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 3150 2746 3206 2748
rect 3230 2746 3286 2748
rect 2990 2694 3036 2746
rect 3036 2694 3046 2746
rect 3070 2694 3100 2746
rect 3100 2694 3112 2746
rect 3112 2694 3126 2746
rect 3150 2694 3164 2746
rect 3164 2694 3176 2746
rect 3176 2694 3206 2746
rect 3230 2694 3240 2746
rect 3240 2694 3286 2746
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 3150 2692 3206 2694
rect 3230 2692 3286 2694
rect 4710 6704 4766 6740
rect 4346 6010 4402 6012
rect 4426 6010 4482 6012
rect 4506 6010 4562 6012
rect 4586 6010 4642 6012
rect 4346 5958 4392 6010
rect 4392 5958 4402 6010
rect 4426 5958 4456 6010
rect 4456 5958 4468 6010
rect 4468 5958 4482 6010
rect 4506 5958 4520 6010
rect 4520 5958 4532 6010
rect 4532 5958 4562 6010
rect 4586 5958 4596 6010
rect 4596 5958 4642 6010
rect 4346 5956 4402 5958
rect 4426 5956 4482 5958
rect 4506 5956 4562 5958
rect 4586 5956 4642 5958
rect 5006 6554 5062 6556
rect 5086 6554 5142 6556
rect 5166 6554 5222 6556
rect 5246 6554 5302 6556
rect 5006 6502 5052 6554
rect 5052 6502 5062 6554
rect 5086 6502 5116 6554
rect 5116 6502 5128 6554
rect 5128 6502 5142 6554
rect 5166 6502 5180 6554
rect 5180 6502 5192 6554
rect 5192 6502 5222 6554
rect 5246 6502 5256 6554
rect 5256 6502 5302 6554
rect 5006 6500 5062 6502
rect 5086 6500 5142 6502
rect 5166 6500 5222 6502
rect 5246 6500 5302 6502
rect 5006 5466 5062 5468
rect 5086 5466 5142 5468
rect 5166 5466 5222 5468
rect 5246 5466 5302 5468
rect 5006 5414 5052 5466
rect 5052 5414 5062 5466
rect 5086 5414 5116 5466
rect 5116 5414 5128 5466
rect 5128 5414 5142 5466
rect 5166 5414 5180 5466
rect 5180 5414 5192 5466
rect 5192 5414 5222 5466
rect 5246 5414 5256 5466
rect 5256 5414 5302 5466
rect 5006 5412 5062 5414
rect 5086 5412 5142 5414
rect 5166 5412 5222 5414
rect 5246 5412 5302 5414
rect 5702 8186 5758 8188
rect 5782 8186 5838 8188
rect 5862 8186 5918 8188
rect 5942 8186 5998 8188
rect 5702 8134 5748 8186
rect 5748 8134 5758 8186
rect 5782 8134 5812 8186
rect 5812 8134 5824 8186
rect 5824 8134 5838 8186
rect 5862 8134 5876 8186
rect 5876 8134 5888 8186
rect 5888 8134 5918 8186
rect 5942 8134 5952 8186
rect 5952 8134 5998 8186
rect 5702 8132 5758 8134
rect 5782 8132 5838 8134
rect 5862 8132 5918 8134
rect 5942 8132 5998 8134
rect 6734 8744 6790 8800
rect 6362 8730 6418 8732
rect 6442 8730 6498 8732
rect 6522 8730 6578 8732
rect 6602 8730 6658 8732
rect 6362 8678 6408 8730
rect 6408 8678 6418 8730
rect 6442 8678 6472 8730
rect 6472 8678 6484 8730
rect 6484 8678 6498 8730
rect 6522 8678 6536 8730
rect 6536 8678 6548 8730
rect 6548 8678 6578 8730
rect 6602 8678 6612 8730
rect 6612 8678 6658 8730
rect 6362 8676 6418 8678
rect 6442 8676 6498 8678
rect 6522 8676 6578 8678
rect 6602 8676 6658 8678
rect 6362 7642 6418 7644
rect 6442 7642 6498 7644
rect 6522 7642 6578 7644
rect 6602 7642 6658 7644
rect 6362 7590 6408 7642
rect 6408 7590 6418 7642
rect 6442 7590 6472 7642
rect 6472 7590 6484 7642
rect 6484 7590 6498 7642
rect 6522 7590 6536 7642
rect 6536 7590 6548 7642
rect 6548 7590 6578 7642
rect 6602 7590 6612 7642
rect 6612 7590 6658 7642
rect 6362 7588 6418 7590
rect 6442 7588 6498 7590
rect 6522 7588 6578 7590
rect 6602 7588 6658 7590
rect 6182 7384 6238 7440
rect 5702 7098 5758 7100
rect 5782 7098 5838 7100
rect 5862 7098 5918 7100
rect 5942 7098 5998 7100
rect 5702 7046 5748 7098
rect 5748 7046 5758 7098
rect 5782 7046 5812 7098
rect 5812 7046 5824 7098
rect 5824 7046 5838 7098
rect 5862 7046 5876 7098
rect 5876 7046 5888 7098
rect 5888 7046 5918 7098
rect 5942 7046 5952 7098
rect 5952 7046 5998 7098
rect 5702 7044 5758 7046
rect 5782 7044 5838 7046
rect 5862 7044 5918 7046
rect 5942 7044 5998 7046
rect 6362 6554 6418 6556
rect 6442 6554 6498 6556
rect 6522 6554 6578 6556
rect 6602 6554 6658 6556
rect 6362 6502 6408 6554
rect 6408 6502 6418 6554
rect 6442 6502 6472 6554
rect 6472 6502 6484 6554
rect 6484 6502 6498 6554
rect 6522 6502 6536 6554
rect 6536 6502 6548 6554
rect 6548 6502 6578 6554
rect 6602 6502 6612 6554
rect 6612 6502 6658 6554
rect 6362 6500 6418 6502
rect 6442 6500 6498 6502
rect 6522 6500 6578 6502
rect 6602 6500 6658 6502
rect 4346 4922 4402 4924
rect 4426 4922 4482 4924
rect 4506 4922 4562 4924
rect 4586 4922 4642 4924
rect 4346 4870 4392 4922
rect 4392 4870 4402 4922
rect 4426 4870 4456 4922
rect 4456 4870 4468 4922
rect 4468 4870 4482 4922
rect 4506 4870 4520 4922
rect 4520 4870 4532 4922
rect 4532 4870 4562 4922
rect 4586 4870 4596 4922
rect 4596 4870 4642 4922
rect 4346 4868 4402 4870
rect 4426 4868 4482 4870
rect 4506 4868 4562 4870
rect 4586 4868 4642 4870
rect 4346 3834 4402 3836
rect 4426 3834 4482 3836
rect 4506 3834 4562 3836
rect 4586 3834 4642 3836
rect 4346 3782 4392 3834
rect 4392 3782 4402 3834
rect 4426 3782 4456 3834
rect 4456 3782 4468 3834
rect 4468 3782 4482 3834
rect 4506 3782 4520 3834
rect 4520 3782 4532 3834
rect 4532 3782 4562 3834
rect 4586 3782 4596 3834
rect 4596 3782 4642 3834
rect 4346 3780 4402 3782
rect 4426 3780 4482 3782
rect 4506 3780 4562 3782
rect 4586 3780 4642 3782
rect 6090 6060 6092 6080
rect 6092 6060 6144 6080
rect 6144 6060 6146 6080
rect 6090 6024 6146 6060
rect 5702 6010 5758 6012
rect 5782 6010 5838 6012
rect 5862 6010 5918 6012
rect 5942 6010 5998 6012
rect 5702 5958 5748 6010
rect 5748 5958 5758 6010
rect 5782 5958 5812 6010
rect 5812 5958 5824 6010
rect 5824 5958 5838 6010
rect 5862 5958 5876 6010
rect 5876 5958 5888 6010
rect 5888 5958 5918 6010
rect 5942 5958 5952 6010
rect 5952 5958 5998 6010
rect 5702 5956 5758 5958
rect 5782 5956 5838 5958
rect 5862 5956 5918 5958
rect 5942 5956 5998 5958
rect 5006 4378 5062 4380
rect 5086 4378 5142 4380
rect 5166 4378 5222 4380
rect 5246 4378 5302 4380
rect 5006 4326 5052 4378
rect 5052 4326 5062 4378
rect 5086 4326 5116 4378
rect 5116 4326 5128 4378
rect 5128 4326 5142 4378
rect 5166 4326 5180 4378
rect 5180 4326 5192 4378
rect 5192 4326 5222 4378
rect 5246 4326 5256 4378
rect 5256 4326 5302 4378
rect 5006 4324 5062 4326
rect 5086 4324 5142 4326
rect 5166 4324 5222 4326
rect 5246 4324 5302 4326
rect 4894 4156 4896 4176
rect 4896 4156 4948 4176
rect 4948 4156 4950 4176
rect 4894 4120 4950 4156
rect 5006 3290 5062 3292
rect 5086 3290 5142 3292
rect 5166 3290 5222 3292
rect 5246 3290 5302 3292
rect 5006 3238 5052 3290
rect 5052 3238 5062 3290
rect 5086 3238 5116 3290
rect 5116 3238 5128 3290
rect 5128 3238 5142 3290
rect 5166 3238 5180 3290
rect 5180 3238 5192 3290
rect 5192 3238 5222 3290
rect 5246 3238 5256 3290
rect 5256 3238 5302 3290
rect 5006 3236 5062 3238
rect 5086 3236 5142 3238
rect 5166 3236 5222 3238
rect 5246 3236 5302 3238
rect 5702 4922 5758 4924
rect 5782 4922 5838 4924
rect 5862 4922 5918 4924
rect 5942 4922 5998 4924
rect 5702 4870 5748 4922
rect 5748 4870 5758 4922
rect 5782 4870 5812 4922
rect 5812 4870 5824 4922
rect 5824 4870 5838 4922
rect 5862 4870 5876 4922
rect 5876 4870 5888 4922
rect 5888 4870 5918 4922
rect 5942 4870 5952 4922
rect 5952 4870 5998 4922
rect 5702 4868 5758 4870
rect 5782 4868 5838 4870
rect 5862 4868 5918 4870
rect 5942 4868 5998 4870
rect 6362 5466 6418 5468
rect 6442 5466 6498 5468
rect 6522 5466 6578 5468
rect 6602 5466 6658 5468
rect 6362 5414 6408 5466
rect 6408 5414 6418 5466
rect 6442 5414 6472 5466
rect 6472 5414 6484 5466
rect 6484 5414 6498 5466
rect 6522 5414 6536 5466
rect 6536 5414 6548 5466
rect 6548 5414 6578 5466
rect 6602 5414 6612 5466
rect 6612 5414 6658 5466
rect 6362 5412 6418 5414
rect 6442 5412 6498 5414
rect 6522 5412 6578 5414
rect 6602 5412 6658 5414
rect 6182 4664 6238 4720
rect 5702 3834 5758 3836
rect 5782 3834 5838 3836
rect 5862 3834 5918 3836
rect 5942 3834 5998 3836
rect 5702 3782 5748 3834
rect 5748 3782 5758 3834
rect 5782 3782 5812 3834
rect 5812 3782 5824 3834
rect 5824 3782 5838 3834
rect 5862 3782 5876 3834
rect 5876 3782 5888 3834
rect 5888 3782 5918 3834
rect 5942 3782 5952 3834
rect 5952 3782 5998 3834
rect 5702 3780 5758 3782
rect 5782 3780 5838 3782
rect 5862 3780 5918 3782
rect 5942 3780 5998 3782
rect 5814 3576 5870 3632
rect 6362 4378 6418 4380
rect 6442 4378 6498 4380
rect 6522 4378 6578 4380
rect 6602 4378 6658 4380
rect 6362 4326 6408 4378
rect 6408 4326 6418 4378
rect 6442 4326 6472 4378
rect 6472 4326 6484 4378
rect 6484 4326 6498 4378
rect 6522 4326 6536 4378
rect 6536 4326 6548 4378
rect 6548 4326 6578 4378
rect 6602 4326 6612 4378
rect 6612 4326 6658 4378
rect 6362 4324 6418 4326
rect 6442 4324 6498 4326
rect 6522 4324 6578 4326
rect 6602 4324 6658 4326
rect 6734 3304 6790 3360
rect 6362 3290 6418 3292
rect 6442 3290 6498 3292
rect 6522 3290 6578 3292
rect 6602 3290 6658 3292
rect 6362 3238 6408 3290
rect 6408 3238 6418 3290
rect 6442 3238 6472 3290
rect 6472 3238 6484 3290
rect 6484 3238 6498 3290
rect 6522 3238 6536 3290
rect 6536 3238 6548 3290
rect 6548 3238 6578 3290
rect 6602 3238 6612 3290
rect 6612 3238 6658 3290
rect 6362 3236 6418 3238
rect 6442 3236 6498 3238
rect 6522 3236 6578 3238
rect 6602 3236 6658 3238
rect 4346 2746 4402 2748
rect 4426 2746 4482 2748
rect 4506 2746 4562 2748
rect 4586 2746 4642 2748
rect 4346 2694 4392 2746
rect 4392 2694 4402 2746
rect 4426 2694 4456 2746
rect 4456 2694 4468 2746
rect 4468 2694 4482 2746
rect 4506 2694 4520 2746
rect 4520 2694 4532 2746
rect 4532 2694 4562 2746
rect 4586 2694 4596 2746
rect 4596 2694 4642 2746
rect 4346 2692 4402 2694
rect 4426 2692 4482 2694
rect 4506 2692 4562 2694
rect 4586 2692 4642 2694
rect 5702 2746 5758 2748
rect 5782 2746 5838 2748
rect 5862 2746 5918 2748
rect 5942 2746 5998 2748
rect 5702 2694 5748 2746
rect 5748 2694 5758 2746
rect 5782 2694 5812 2746
rect 5812 2694 5824 2746
rect 5824 2694 5838 2746
rect 5862 2694 5876 2746
rect 5876 2694 5888 2746
rect 5888 2694 5918 2746
rect 5942 2694 5952 2746
rect 5952 2694 5998 2746
rect 5702 2692 5758 2694
rect 5782 2692 5838 2694
rect 5862 2692 5918 2694
rect 5942 2692 5998 2694
rect 3650 2202 3706 2204
rect 3730 2202 3786 2204
rect 3810 2202 3866 2204
rect 3890 2202 3946 2204
rect 3650 2150 3696 2202
rect 3696 2150 3706 2202
rect 3730 2150 3760 2202
rect 3760 2150 3772 2202
rect 3772 2150 3786 2202
rect 3810 2150 3824 2202
rect 3824 2150 3836 2202
rect 3836 2150 3866 2202
rect 3890 2150 3900 2202
rect 3900 2150 3946 2202
rect 3650 2148 3706 2150
rect 3730 2148 3786 2150
rect 3810 2148 3866 2150
rect 3890 2148 3946 2150
rect 5006 2202 5062 2204
rect 5086 2202 5142 2204
rect 5166 2202 5222 2204
rect 5246 2202 5302 2204
rect 5006 2150 5052 2202
rect 5052 2150 5062 2202
rect 5086 2150 5116 2202
rect 5116 2150 5128 2202
rect 5128 2150 5142 2202
rect 5166 2150 5180 2202
rect 5180 2150 5192 2202
rect 5192 2150 5222 2202
rect 5246 2150 5256 2202
rect 5256 2150 5302 2202
rect 5006 2148 5062 2150
rect 5086 2148 5142 2150
rect 5166 2148 5222 2150
rect 5246 2148 5302 2150
rect 5538 1944 5594 2000
rect 2778 1400 2834 1456
rect 6362 2202 6418 2204
rect 6442 2202 6498 2204
rect 6522 2202 6578 2204
rect 6602 2202 6658 2204
rect 6362 2150 6408 2202
rect 6408 2150 6418 2202
rect 6442 2150 6472 2202
rect 6472 2150 6484 2202
rect 6484 2150 6498 2202
rect 6522 2150 6536 2202
rect 6536 2150 6548 2202
rect 6548 2150 6578 2202
rect 6602 2150 6612 2202
rect 6612 2150 6658 2202
rect 6362 2148 6418 2150
rect 6442 2148 6498 2150
rect 6522 2148 6578 2150
rect 6602 2148 6658 2150
rect 6182 584 6238 640
<< metal3 >>
rect 6361 11522 6427 11525
rect 6901 11522 7701 11552
rect 6361 11520 7701 11522
rect 6361 11464 6366 11520
rect 6422 11464 7701 11520
rect 6361 11462 7701 11464
rect 6361 11459 6427 11462
rect 6901 11432 7701 11462
rect 0 10978 800 11008
rect 933 10978 999 10981
rect 0 10976 999 10978
rect 0 10920 938 10976
rect 994 10920 999 10976
rect 0 10918 999 10920
rect 0 10888 800 10918
rect 933 10915 999 10918
rect 1624 10368 1940 10369
rect 1624 10304 1630 10368
rect 1694 10304 1710 10368
rect 1774 10304 1790 10368
rect 1854 10304 1870 10368
rect 1934 10304 1940 10368
rect 1624 10303 1940 10304
rect 2980 10368 3296 10369
rect 2980 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3146 10368
rect 3210 10304 3226 10368
rect 3290 10304 3296 10368
rect 2980 10303 3296 10304
rect 4336 10368 4652 10369
rect 4336 10304 4342 10368
rect 4406 10304 4422 10368
rect 4486 10304 4502 10368
rect 4566 10304 4582 10368
rect 4646 10304 4652 10368
rect 4336 10303 4652 10304
rect 5692 10368 6008 10369
rect 5692 10304 5698 10368
rect 5762 10304 5778 10368
rect 5842 10304 5858 10368
rect 5922 10304 5938 10368
rect 6002 10304 6008 10368
rect 5692 10303 6008 10304
rect 5349 10162 5415 10165
rect 6901 10162 7701 10192
rect 5349 10160 7701 10162
rect 5349 10104 5354 10160
rect 5410 10104 7701 10160
rect 5349 10102 7701 10104
rect 5349 10099 5415 10102
rect 6901 10072 7701 10102
rect 2284 9824 2600 9825
rect 2284 9760 2290 9824
rect 2354 9760 2370 9824
rect 2434 9760 2450 9824
rect 2514 9760 2530 9824
rect 2594 9760 2600 9824
rect 2284 9759 2600 9760
rect 3640 9824 3956 9825
rect 3640 9760 3646 9824
rect 3710 9760 3726 9824
rect 3790 9760 3806 9824
rect 3870 9760 3886 9824
rect 3950 9760 3956 9824
rect 3640 9759 3956 9760
rect 4996 9824 5312 9825
rect 4996 9760 5002 9824
rect 5066 9760 5082 9824
rect 5146 9760 5162 9824
rect 5226 9760 5242 9824
rect 5306 9760 5312 9824
rect 4996 9759 5312 9760
rect 6352 9824 6668 9825
rect 6352 9760 6358 9824
rect 6422 9760 6438 9824
rect 6502 9760 6518 9824
rect 6582 9760 6598 9824
rect 6662 9760 6668 9824
rect 6352 9759 6668 9760
rect 1624 9280 1940 9281
rect 1624 9216 1630 9280
rect 1694 9216 1710 9280
rect 1774 9216 1790 9280
rect 1854 9216 1870 9280
rect 1934 9216 1940 9280
rect 1624 9215 1940 9216
rect 2980 9280 3296 9281
rect 2980 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3146 9280
rect 3210 9216 3226 9280
rect 3290 9216 3296 9280
rect 2980 9215 3296 9216
rect 4336 9280 4652 9281
rect 4336 9216 4342 9280
rect 4406 9216 4422 9280
rect 4486 9216 4502 9280
rect 4566 9216 4582 9280
rect 4646 9216 4652 9280
rect 4336 9215 4652 9216
rect 5692 9280 6008 9281
rect 5692 9216 5698 9280
rect 5762 9216 5778 9280
rect 5842 9216 5858 9280
rect 5922 9216 5938 9280
rect 6002 9216 6008 9280
rect 5692 9215 6008 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 6729 8802 6795 8805
rect 6901 8802 7701 8832
rect 6729 8800 7701 8802
rect 6729 8744 6734 8800
rect 6790 8744 7701 8800
rect 6729 8742 7701 8744
rect 6729 8739 6795 8742
rect 2284 8736 2600 8737
rect 2284 8672 2290 8736
rect 2354 8672 2370 8736
rect 2434 8672 2450 8736
rect 2514 8672 2530 8736
rect 2594 8672 2600 8736
rect 2284 8671 2600 8672
rect 3640 8736 3956 8737
rect 3640 8672 3646 8736
rect 3710 8672 3726 8736
rect 3790 8672 3806 8736
rect 3870 8672 3886 8736
rect 3950 8672 3956 8736
rect 3640 8671 3956 8672
rect 4996 8736 5312 8737
rect 4996 8672 5002 8736
rect 5066 8672 5082 8736
rect 5146 8672 5162 8736
rect 5226 8672 5242 8736
rect 5306 8672 5312 8736
rect 4996 8671 5312 8672
rect 6352 8736 6668 8737
rect 6352 8672 6358 8736
rect 6422 8672 6438 8736
rect 6502 8672 6518 8736
rect 6582 8672 6598 8736
rect 6662 8672 6668 8736
rect 6901 8712 7701 8742
rect 6352 8671 6668 8672
rect 1624 8192 1940 8193
rect 1624 8128 1630 8192
rect 1694 8128 1710 8192
rect 1774 8128 1790 8192
rect 1854 8128 1870 8192
rect 1934 8128 1940 8192
rect 1624 8127 1940 8128
rect 2980 8192 3296 8193
rect 2980 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3146 8192
rect 3210 8128 3226 8192
rect 3290 8128 3296 8192
rect 2980 8127 3296 8128
rect 4336 8192 4652 8193
rect 4336 8128 4342 8192
rect 4406 8128 4422 8192
rect 4486 8128 4502 8192
rect 4566 8128 4582 8192
rect 4646 8128 4652 8192
rect 4336 8127 4652 8128
rect 5692 8192 6008 8193
rect 5692 8128 5698 8192
rect 5762 8128 5778 8192
rect 5842 8128 5858 8192
rect 5922 8128 5938 8192
rect 6002 8128 6008 8192
rect 5692 8127 6008 8128
rect 2284 7648 2600 7649
rect 2284 7584 2290 7648
rect 2354 7584 2370 7648
rect 2434 7584 2450 7648
rect 2514 7584 2530 7648
rect 2594 7584 2600 7648
rect 2284 7583 2600 7584
rect 3640 7648 3956 7649
rect 3640 7584 3646 7648
rect 3710 7584 3726 7648
rect 3790 7584 3806 7648
rect 3870 7584 3886 7648
rect 3950 7584 3956 7648
rect 3640 7583 3956 7584
rect 4996 7648 5312 7649
rect 4996 7584 5002 7648
rect 5066 7584 5082 7648
rect 5146 7584 5162 7648
rect 5226 7584 5242 7648
rect 5306 7584 5312 7648
rect 4996 7583 5312 7584
rect 6352 7648 6668 7649
rect 6352 7584 6358 7648
rect 6422 7584 6438 7648
rect 6502 7584 6518 7648
rect 6582 7584 6598 7648
rect 6662 7584 6668 7648
rect 6352 7583 6668 7584
rect 6177 7442 6243 7445
rect 6901 7442 7701 7472
rect 6177 7440 7701 7442
rect 6177 7384 6182 7440
rect 6238 7384 7701 7440
rect 6177 7382 7701 7384
rect 6177 7379 6243 7382
rect 6901 7352 7701 7382
rect 0 7170 800 7200
rect 0 7080 858 7170
rect 798 7034 858 7080
rect 1624 7104 1940 7105
rect 1624 7040 1630 7104
rect 1694 7040 1710 7104
rect 1774 7040 1790 7104
rect 1854 7040 1870 7104
rect 1934 7040 1940 7104
rect 1624 7039 1940 7040
rect 2980 7104 3296 7105
rect 2980 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3146 7104
rect 3210 7040 3226 7104
rect 3290 7040 3296 7104
rect 2980 7039 3296 7040
rect 4336 7104 4652 7105
rect 4336 7040 4342 7104
rect 4406 7040 4422 7104
rect 4486 7040 4502 7104
rect 4566 7040 4582 7104
rect 4646 7040 4652 7104
rect 4336 7039 4652 7040
rect 5692 7104 6008 7105
rect 5692 7040 5698 7104
rect 5762 7040 5778 7104
rect 5842 7040 5858 7104
rect 5922 7040 5938 7104
rect 6002 7040 6008 7104
rect 5692 7039 6008 7040
rect 1393 7034 1459 7037
rect 798 7032 1459 7034
rect 798 6976 1398 7032
rect 1454 6976 1459 7032
rect 798 6974 1459 6976
rect 1393 6971 1459 6974
rect 2681 6898 2747 6901
rect 4245 6898 4311 6901
rect 2681 6896 4311 6898
rect 2681 6840 2686 6896
rect 2742 6840 4250 6896
rect 4306 6840 4311 6896
rect 2681 6838 4311 6840
rect 2681 6835 2747 6838
rect 4245 6835 4311 6838
rect 2221 6762 2287 6765
rect 4705 6762 4771 6765
rect 2221 6760 4771 6762
rect 2221 6704 2226 6760
rect 2282 6704 4710 6760
rect 4766 6704 4771 6760
rect 2221 6702 4771 6704
rect 2221 6699 2287 6702
rect 4705 6699 4771 6702
rect 2284 6560 2600 6561
rect 2284 6496 2290 6560
rect 2354 6496 2370 6560
rect 2434 6496 2450 6560
rect 2514 6496 2530 6560
rect 2594 6496 2600 6560
rect 2284 6495 2600 6496
rect 3640 6560 3956 6561
rect 3640 6496 3646 6560
rect 3710 6496 3726 6560
rect 3790 6496 3806 6560
rect 3870 6496 3886 6560
rect 3950 6496 3956 6560
rect 3640 6495 3956 6496
rect 4996 6560 5312 6561
rect 4996 6496 5002 6560
rect 5066 6496 5082 6560
rect 5146 6496 5162 6560
rect 5226 6496 5242 6560
rect 5306 6496 5312 6560
rect 4996 6495 5312 6496
rect 6352 6560 6668 6561
rect 6352 6496 6358 6560
rect 6422 6496 6438 6560
rect 6502 6496 6518 6560
rect 6582 6496 6598 6560
rect 6662 6496 6668 6560
rect 6352 6495 6668 6496
rect 6085 6082 6151 6085
rect 6901 6082 7701 6112
rect 6085 6080 7701 6082
rect 6085 6024 6090 6080
rect 6146 6024 7701 6080
rect 6085 6022 7701 6024
rect 6085 6019 6151 6022
rect 1624 6016 1940 6017
rect 1624 5952 1630 6016
rect 1694 5952 1710 6016
rect 1774 5952 1790 6016
rect 1854 5952 1870 6016
rect 1934 5952 1940 6016
rect 1624 5951 1940 5952
rect 2980 6016 3296 6017
rect 2980 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3146 6016
rect 3210 5952 3226 6016
rect 3290 5952 3296 6016
rect 2980 5951 3296 5952
rect 4336 6016 4652 6017
rect 4336 5952 4342 6016
rect 4406 5952 4422 6016
rect 4486 5952 4502 6016
rect 4566 5952 4582 6016
rect 4646 5952 4652 6016
rect 4336 5951 4652 5952
rect 5692 6016 6008 6017
rect 5692 5952 5698 6016
rect 5762 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5938 6016
rect 6002 5952 6008 6016
rect 6901 5992 7701 6022
rect 5692 5951 6008 5952
rect 1393 5536 1459 5541
rect 1393 5480 1398 5536
rect 1454 5480 1459 5536
rect 1393 5475 1459 5480
rect 0 5266 800 5296
rect 1396 5266 1456 5475
rect 2284 5472 2600 5473
rect 2284 5408 2290 5472
rect 2354 5408 2370 5472
rect 2434 5408 2450 5472
rect 2514 5408 2530 5472
rect 2594 5408 2600 5472
rect 2284 5407 2600 5408
rect 3640 5472 3956 5473
rect 3640 5408 3646 5472
rect 3710 5408 3726 5472
rect 3790 5408 3806 5472
rect 3870 5408 3886 5472
rect 3950 5408 3956 5472
rect 3640 5407 3956 5408
rect 4996 5472 5312 5473
rect 4996 5408 5002 5472
rect 5066 5408 5082 5472
rect 5146 5408 5162 5472
rect 5226 5408 5242 5472
rect 5306 5408 5312 5472
rect 4996 5407 5312 5408
rect 6352 5472 6668 5473
rect 6352 5408 6358 5472
rect 6422 5408 6438 5472
rect 6502 5408 6518 5472
rect 6582 5408 6598 5472
rect 6662 5408 6668 5472
rect 6352 5407 6668 5408
rect 0 5206 1456 5266
rect 0 5176 800 5206
rect 1624 4928 1940 4929
rect 1624 4864 1630 4928
rect 1694 4864 1710 4928
rect 1774 4864 1790 4928
rect 1854 4864 1870 4928
rect 1934 4864 1940 4928
rect 1624 4863 1940 4864
rect 2980 4928 3296 4929
rect 2980 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3146 4928
rect 3210 4864 3226 4928
rect 3290 4864 3296 4928
rect 2980 4863 3296 4864
rect 4336 4928 4652 4929
rect 4336 4864 4342 4928
rect 4406 4864 4422 4928
rect 4486 4864 4502 4928
rect 4566 4864 4582 4928
rect 4646 4864 4652 4928
rect 4336 4863 4652 4864
rect 5692 4928 6008 4929
rect 5692 4864 5698 4928
rect 5762 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5938 4928
rect 6002 4864 6008 4928
rect 5692 4863 6008 4864
rect 2681 4722 2747 4725
rect 2957 4722 3023 4725
rect 2681 4720 3023 4722
rect 2681 4664 2686 4720
rect 2742 4664 2962 4720
rect 3018 4664 3023 4720
rect 2681 4662 3023 4664
rect 2681 4659 2747 4662
rect 2957 4659 3023 4662
rect 6177 4722 6243 4725
rect 6901 4722 7701 4752
rect 6177 4720 7701 4722
rect 6177 4664 6182 4720
rect 6238 4664 7701 4720
rect 6177 4662 7701 4664
rect 6177 4659 6243 4662
rect 6901 4632 7701 4662
rect 2284 4384 2600 4385
rect 2284 4320 2290 4384
rect 2354 4320 2370 4384
rect 2434 4320 2450 4384
rect 2514 4320 2530 4384
rect 2594 4320 2600 4384
rect 2284 4319 2600 4320
rect 3640 4384 3956 4385
rect 3640 4320 3646 4384
rect 3710 4320 3726 4384
rect 3790 4320 3806 4384
rect 3870 4320 3886 4384
rect 3950 4320 3956 4384
rect 3640 4319 3956 4320
rect 4996 4384 5312 4385
rect 4996 4320 5002 4384
rect 5066 4320 5082 4384
rect 5146 4320 5162 4384
rect 5226 4320 5242 4384
rect 5306 4320 5312 4384
rect 4996 4319 5312 4320
rect 6352 4384 6668 4385
rect 6352 4320 6358 4384
rect 6422 4320 6438 4384
rect 6502 4320 6518 4384
rect 6582 4320 6598 4384
rect 6662 4320 6668 4384
rect 6352 4319 6668 4320
rect 2957 4178 3023 4181
rect 4889 4178 4955 4181
rect 2957 4176 4955 4178
rect 2957 4120 2962 4176
rect 3018 4120 4894 4176
rect 4950 4120 4955 4176
rect 2957 4118 4955 4120
rect 2957 4115 3023 4118
rect 4889 4115 4955 4118
rect 1624 3840 1940 3841
rect 1624 3776 1630 3840
rect 1694 3776 1710 3840
rect 1774 3776 1790 3840
rect 1854 3776 1870 3840
rect 1934 3776 1940 3840
rect 1624 3775 1940 3776
rect 2980 3840 3296 3841
rect 2980 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3146 3840
rect 3210 3776 3226 3840
rect 3290 3776 3296 3840
rect 2980 3775 3296 3776
rect 4336 3840 4652 3841
rect 4336 3776 4342 3840
rect 4406 3776 4422 3840
rect 4486 3776 4502 3840
rect 4566 3776 4582 3840
rect 4646 3776 4652 3840
rect 4336 3775 4652 3776
rect 5692 3840 6008 3841
rect 5692 3776 5698 3840
rect 5762 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5938 3840
rect 6002 3776 6008 3840
rect 5692 3775 6008 3776
rect 2681 3634 2747 3637
rect 5809 3634 5875 3637
rect 2681 3632 5875 3634
rect 2681 3576 2686 3632
rect 2742 3576 5814 3632
rect 5870 3576 5875 3632
rect 2681 3574 5875 3576
rect 2681 3571 2747 3574
rect 5809 3571 5875 3574
rect 0 3362 800 3392
rect 933 3362 999 3365
rect 0 3360 999 3362
rect 0 3304 938 3360
rect 994 3304 999 3360
rect 0 3302 999 3304
rect 0 3272 800 3302
rect 933 3299 999 3302
rect 6729 3362 6795 3365
rect 6901 3362 7701 3392
rect 6729 3360 7701 3362
rect 6729 3304 6734 3360
rect 6790 3304 7701 3360
rect 6729 3302 7701 3304
rect 6729 3299 6795 3302
rect 2284 3296 2600 3297
rect 2284 3232 2290 3296
rect 2354 3232 2370 3296
rect 2434 3232 2450 3296
rect 2514 3232 2530 3296
rect 2594 3232 2600 3296
rect 2284 3231 2600 3232
rect 3640 3296 3956 3297
rect 3640 3232 3646 3296
rect 3710 3232 3726 3296
rect 3790 3232 3806 3296
rect 3870 3232 3886 3296
rect 3950 3232 3956 3296
rect 3640 3231 3956 3232
rect 4996 3296 5312 3297
rect 4996 3232 5002 3296
rect 5066 3232 5082 3296
rect 5146 3232 5162 3296
rect 5226 3232 5242 3296
rect 5306 3232 5312 3296
rect 4996 3231 5312 3232
rect 6352 3296 6668 3297
rect 6352 3232 6358 3296
rect 6422 3232 6438 3296
rect 6502 3232 6518 3296
rect 6582 3232 6598 3296
rect 6662 3232 6668 3296
rect 6901 3272 7701 3302
rect 6352 3231 6668 3232
rect 1624 2752 1940 2753
rect 1624 2688 1630 2752
rect 1694 2688 1710 2752
rect 1774 2688 1790 2752
rect 1854 2688 1870 2752
rect 1934 2688 1940 2752
rect 1624 2687 1940 2688
rect 2980 2752 3296 2753
rect 2980 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3146 2752
rect 3210 2688 3226 2752
rect 3290 2688 3296 2752
rect 2980 2687 3296 2688
rect 4336 2752 4652 2753
rect 4336 2688 4342 2752
rect 4406 2688 4422 2752
rect 4486 2688 4502 2752
rect 4566 2688 4582 2752
rect 4646 2688 4652 2752
rect 4336 2687 4652 2688
rect 5692 2752 6008 2753
rect 5692 2688 5698 2752
rect 5762 2688 5778 2752
rect 5842 2688 5858 2752
rect 5922 2688 5938 2752
rect 6002 2688 6008 2752
rect 5692 2687 6008 2688
rect 2284 2208 2600 2209
rect 2284 2144 2290 2208
rect 2354 2144 2370 2208
rect 2434 2144 2450 2208
rect 2514 2144 2530 2208
rect 2594 2144 2600 2208
rect 2284 2143 2600 2144
rect 3640 2208 3956 2209
rect 3640 2144 3646 2208
rect 3710 2144 3726 2208
rect 3790 2144 3806 2208
rect 3870 2144 3886 2208
rect 3950 2144 3956 2208
rect 3640 2143 3956 2144
rect 4996 2208 5312 2209
rect 4996 2144 5002 2208
rect 5066 2144 5082 2208
rect 5146 2144 5162 2208
rect 5226 2144 5242 2208
rect 5306 2144 5312 2208
rect 4996 2143 5312 2144
rect 6352 2208 6668 2209
rect 6352 2144 6358 2208
rect 6422 2144 6438 2208
rect 6502 2144 6518 2208
rect 6582 2144 6598 2208
rect 6662 2144 6668 2208
rect 6352 2143 6668 2144
rect 5533 2002 5599 2005
rect 6901 2002 7701 2032
rect 5533 2000 7701 2002
rect 5533 1944 5538 2000
rect 5594 1944 7701 2000
rect 5533 1942 7701 1944
rect 5533 1939 5599 1942
rect 6901 1912 7701 1942
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 6177 642 6243 645
rect 6901 642 7701 672
rect 6177 640 7701 642
rect 6177 584 6182 640
rect 6238 584 7701 640
rect 6177 582 7701 584
rect 6177 579 6243 582
rect 6901 552 7701 582
<< via3 >>
rect 1630 10364 1694 10368
rect 1630 10308 1634 10364
rect 1634 10308 1690 10364
rect 1690 10308 1694 10364
rect 1630 10304 1694 10308
rect 1710 10364 1774 10368
rect 1710 10308 1714 10364
rect 1714 10308 1770 10364
rect 1770 10308 1774 10364
rect 1710 10304 1774 10308
rect 1790 10364 1854 10368
rect 1790 10308 1794 10364
rect 1794 10308 1850 10364
rect 1850 10308 1854 10364
rect 1790 10304 1854 10308
rect 1870 10364 1934 10368
rect 1870 10308 1874 10364
rect 1874 10308 1930 10364
rect 1930 10308 1934 10364
rect 1870 10304 1934 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 3146 10364 3210 10368
rect 3146 10308 3150 10364
rect 3150 10308 3206 10364
rect 3206 10308 3210 10364
rect 3146 10304 3210 10308
rect 3226 10364 3290 10368
rect 3226 10308 3230 10364
rect 3230 10308 3286 10364
rect 3286 10308 3290 10364
rect 3226 10304 3290 10308
rect 4342 10364 4406 10368
rect 4342 10308 4346 10364
rect 4346 10308 4402 10364
rect 4402 10308 4406 10364
rect 4342 10304 4406 10308
rect 4422 10364 4486 10368
rect 4422 10308 4426 10364
rect 4426 10308 4482 10364
rect 4482 10308 4486 10364
rect 4422 10304 4486 10308
rect 4502 10364 4566 10368
rect 4502 10308 4506 10364
rect 4506 10308 4562 10364
rect 4562 10308 4566 10364
rect 4502 10304 4566 10308
rect 4582 10364 4646 10368
rect 4582 10308 4586 10364
rect 4586 10308 4642 10364
rect 4642 10308 4646 10364
rect 4582 10304 4646 10308
rect 5698 10364 5762 10368
rect 5698 10308 5702 10364
rect 5702 10308 5758 10364
rect 5758 10308 5762 10364
rect 5698 10304 5762 10308
rect 5778 10364 5842 10368
rect 5778 10308 5782 10364
rect 5782 10308 5838 10364
rect 5838 10308 5842 10364
rect 5778 10304 5842 10308
rect 5858 10364 5922 10368
rect 5858 10308 5862 10364
rect 5862 10308 5918 10364
rect 5918 10308 5922 10364
rect 5858 10304 5922 10308
rect 5938 10364 6002 10368
rect 5938 10308 5942 10364
rect 5942 10308 5998 10364
rect 5998 10308 6002 10364
rect 5938 10304 6002 10308
rect 2290 9820 2354 9824
rect 2290 9764 2294 9820
rect 2294 9764 2350 9820
rect 2350 9764 2354 9820
rect 2290 9760 2354 9764
rect 2370 9820 2434 9824
rect 2370 9764 2374 9820
rect 2374 9764 2430 9820
rect 2430 9764 2434 9820
rect 2370 9760 2434 9764
rect 2450 9820 2514 9824
rect 2450 9764 2454 9820
rect 2454 9764 2510 9820
rect 2510 9764 2514 9820
rect 2450 9760 2514 9764
rect 2530 9820 2594 9824
rect 2530 9764 2534 9820
rect 2534 9764 2590 9820
rect 2590 9764 2594 9820
rect 2530 9760 2594 9764
rect 3646 9820 3710 9824
rect 3646 9764 3650 9820
rect 3650 9764 3706 9820
rect 3706 9764 3710 9820
rect 3646 9760 3710 9764
rect 3726 9820 3790 9824
rect 3726 9764 3730 9820
rect 3730 9764 3786 9820
rect 3786 9764 3790 9820
rect 3726 9760 3790 9764
rect 3806 9820 3870 9824
rect 3806 9764 3810 9820
rect 3810 9764 3866 9820
rect 3866 9764 3870 9820
rect 3806 9760 3870 9764
rect 3886 9820 3950 9824
rect 3886 9764 3890 9820
rect 3890 9764 3946 9820
rect 3946 9764 3950 9820
rect 3886 9760 3950 9764
rect 5002 9820 5066 9824
rect 5002 9764 5006 9820
rect 5006 9764 5062 9820
rect 5062 9764 5066 9820
rect 5002 9760 5066 9764
rect 5082 9820 5146 9824
rect 5082 9764 5086 9820
rect 5086 9764 5142 9820
rect 5142 9764 5146 9820
rect 5082 9760 5146 9764
rect 5162 9820 5226 9824
rect 5162 9764 5166 9820
rect 5166 9764 5222 9820
rect 5222 9764 5226 9820
rect 5162 9760 5226 9764
rect 5242 9820 5306 9824
rect 5242 9764 5246 9820
rect 5246 9764 5302 9820
rect 5302 9764 5306 9820
rect 5242 9760 5306 9764
rect 6358 9820 6422 9824
rect 6358 9764 6362 9820
rect 6362 9764 6418 9820
rect 6418 9764 6422 9820
rect 6358 9760 6422 9764
rect 6438 9820 6502 9824
rect 6438 9764 6442 9820
rect 6442 9764 6498 9820
rect 6498 9764 6502 9820
rect 6438 9760 6502 9764
rect 6518 9820 6582 9824
rect 6518 9764 6522 9820
rect 6522 9764 6578 9820
rect 6578 9764 6582 9820
rect 6518 9760 6582 9764
rect 6598 9820 6662 9824
rect 6598 9764 6602 9820
rect 6602 9764 6658 9820
rect 6658 9764 6662 9820
rect 6598 9760 6662 9764
rect 1630 9276 1694 9280
rect 1630 9220 1634 9276
rect 1634 9220 1690 9276
rect 1690 9220 1694 9276
rect 1630 9216 1694 9220
rect 1710 9276 1774 9280
rect 1710 9220 1714 9276
rect 1714 9220 1770 9276
rect 1770 9220 1774 9276
rect 1710 9216 1774 9220
rect 1790 9276 1854 9280
rect 1790 9220 1794 9276
rect 1794 9220 1850 9276
rect 1850 9220 1854 9276
rect 1790 9216 1854 9220
rect 1870 9276 1934 9280
rect 1870 9220 1874 9276
rect 1874 9220 1930 9276
rect 1930 9220 1934 9276
rect 1870 9216 1934 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 3146 9276 3210 9280
rect 3146 9220 3150 9276
rect 3150 9220 3206 9276
rect 3206 9220 3210 9276
rect 3146 9216 3210 9220
rect 3226 9276 3290 9280
rect 3226 9220 3230 9276
rect 3230 9220 3286 9276
rect 3286 9220 3290 9276
rect 3226 9216 3290 9220
rect 4342 9276 4406 9280
rect 4342 9220 4346 9276
rect 4346 9220 4402 9276
rect 4402 9220 4406 9276
rect 4342 9216 4406 9220
rect 4422 9276 4486 9280
rect 4422 9220 4426 9276
rect 4426 9220 4482 9276
rect 4482 9220 4486 9276
rect 4422 9216 4486 9220
rect 4502 9276 4566 9280
rect 4502 9220 4506 9276
rect 4506 9220 4562 9276
rect 4562 9220 4566 9276
rect 4502 9216 4566 9220
rect 4582 9276 4646 9280
rect 4582 9220 4586 9276
rect 4586 9220 4642 9276
rect 4642 9220 4646 9276
rect 4582 9216 4646 9220
rect 5698 9276 5762 9280
rect 5698 9220 5702 9276
rect 5702 9220 5758 9276
rect 5758 9220 5762 9276
rect 5698 9216 5762 9220
rect 5778 9276 5842 9280
rect 5778 9220 5782 9276
rect 5782 9220 5838 9276
rect 5838 9220 5842 9276
rect 5778 9216 5842 9220
rect 5858 9276 5922 9280
rect 5858 9220 5862 9276
rect 5862 9220 5918 9276
rect 5918 9220 5922 9276
rect 5858 9216 5922 9220
rect 5938 9276 6002 9280
rect 5938 9220 5942 9276
rect 5942 9220 5998 9276
rect 5998 9220 6002 9276
rect 5938 9216 6002 9220
rect 2290 8732 2354 8736
rect 2290 8676 2294 8732
rect 2294 8676 2350 8732
rect 2350 8676 2354 8732
rect 2290 8672 2354 8676
rect 2370 8732 2434 8736
rect 2370 8676 2374 8732
rect 2374 8676 2430 8732
rect 2430 8676 2434 8732
rect 2370 8672 2434 8676
rect 2450 8732 2514 8736
rect 2450 8676 2454 8732
rect 2454 8676 2510 8732
rect 2510 8676 2514 8732
rect 2450 8672 2514 8676
rect 2530 8732 2594 8736
rect 2530 8676 2534 8732
rect 2534 8676 2590 8732
rect 2590 8676 2594 8732
rect 2530 8672 2594 8676
rect 3646 8732 3710 8736
rect 3646 8676 3650 8732
rect 3650 8676 3706 8732
rect 3706 8676 3710 8732
rect 3646 8672 3710 8676
rect 3726 8732 3790 8736
rect 3726 8676 3730 8732
rect 3730 8676 3786 8732
rect 3786 8676 3790 8732
rect 3726 8672 3790 8676
rect 3806 8732 3870 8736
rect 3806 8676 3810 8732
rect 3810 8676 3866 8732
rect 3866 8676 3870 8732
rect 3806 8672 3870 8676
rect 3886 8732 3950 8736
rect 3886 8676 3890 8732
rect 3890 8676 3946 8732
rect 3946 8676 3950 8732
rect 3886 8672 3950 8676
rect 5002 8732 5066 8736
rect 5002 8676 5006 8732
rect 5006 8676 5062 8732
rect 5062 8676 5066 8732
rect 5002 8672 5066 8676
rect 5082 8732 5146 8736
rect 5082 8676 5086 8732
rect 5086 8676 5142 8732
rect 5142 8676 5146 8732
rect 5082 8672 5146 8676
rect 5162 8732 5226 8736
rect 5162 8676 5166 8732
rect 5166 8676 5222 8732
rect 5222 8676 5226 8732
rect 5162 8672 5226 8676
rect 5242 8732 5306 8736
rect 5242 8676 5246 8732
rect 5246 8676 5302 8732
rect 5302 8676 5306 8732
rect 5242 8672 5306 8676
rect 6358 8732 6422 8736
rect 6358 8676 6362 8732
rect 6362 8676 6418 8732
rect 6418 8676 6422 8732
rect 6358 8672 6422 8676
rect 6438 8732 6502 8736
rect 6438 8676 6442 8732
rect 6442 8676 6498 8732
rect 6498 8676 6502 8732
rect 6438 8672 6502 8676
rect 6518 8732 6582 8736
rect 6518 8676 6522 8732
rect 6522 8676 6578 8732
rect 6578 8676 6582 8732
rect 6518 8672 6582 8676
rect 6598 8732 6662 8736
rect 6598 8676 6602 8732
rect 6602 8676 6658 8732
rect 6658 8676 6662 8732
rect 6598 8672 6662 8676
rect 1630 8188 1694 8192
rect 1630 8132 1634 8188
rect 1634 8132 1690 8188
rect 1690 8132 1694 8188
rect 1630 8128 1694 8132
rect 1710 8188 1774 8192
rect 1710 8132 1714 8188
rect 1714 8132 1770 8188
rect 1770 8132 1774 8188
rect 1710 8128 1774 8132
rect 1790 8188 1854 8192
rect 1790 8132 1794 8188
rect 1794 8132 1850 8188
rect 1850 8132 1854 8188
rect 1790 8128 1854 8132
rect 1870 8188 1934 8192
rect 1870 8132 1874 8188
rect 1874 8132 1930 8188
rect 1930 8132 1934 8188
rect 1870 8128 1934 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 3146 8188 3210 8192
rect 3146 8132 3150 8188
rect 3150 8132 3206 8188
rect 3206 8132 3210 8188
rect 3146 8128 3210 8132
rect 3226 8188 3290 8192
rect 3226 8132 3230 8188
rect 3230 8132 3286 8188
rect 3286 8132 3290 8188
rect 3226 8128 3290 8132
rect 4342 8188 4406 8192
rect 4342 8132 4346 8188
rect 4346 8132 4402 8188
rect 4402 8132 4406 8188
rect 4342 8128 4406 8132
rect 4422 8188 4486 8192
rect 4422 8132 4426 8188
rect 4426 8132 4482 8188
rect 4482 8132 4486 8188
rect 4422 8128 4486 8132
rect 4502 8188 4566 8192
rect 4502 8132 4506 8188
rect 4506 8132 4562 8188
rect 4562 8132 4566 8188
rect 4502 8128 4566 8132
rect 4582 8188 4646 8192
rect 4582 8132 4586 8188
rect 4586 8132 4642 8188
rect 4642 8132 4646 8188
rect 4582 8128 4646 8132
rect 5698 8188 5762 8192
rect 5698 8132 5702 8188
rect 5702 8132 5758 8188
rect 5758 8132 5762 8188
rect 5698 8128 5762 8132
rect 5778 8188 5842 8192
rect 5778 8132 5782 8188
rect 5782 8132 5838 8188
rect 5838 8132 5842 8188
rect 5778 8128 5842 8132
rect 5858 8188 5922 8192
rect 5858 8132 5862 8188
rect 5862 8132 5918 8188
rect 5918 8132 5922 8188
rect 5858 8128 5922 8132
rect 5938 8188 6002 8192
rect 5938 8132 5942 8188
rect 5942 8132 5998 8188
rect 5998 8132 6002 8188
rect 5938 8128 6002 8132
rect 2290 7644 2354 7648
rect 2290 7588 2294 7644
rect 2294 7588 2350 7644
rect 2350 7588 2354 7644
rect 2290 7584 2354 7588
rect 2370 7644 2434 7648
rect 2370 7588 2374 7644
rect 2374 7588 2430 7644
rect 2430 7588 2434 7644
rect 2370 7584 2434 7588
rect 2450 7644 2514 7648
rect 2450 7588 2454 7644
rect 2454 7588 2510 7644
rect 2510 7588 2514 7644
rect 2450 7584 2514 7588
rect 2530 7644 2594 7648
rect 2530 7588 2534 7644
rect 2534 7588 2590 7644
rect 2590 7588 2594 7644
rect 2530 7584 2594 7588
rect 3646 7644 3710 7648
rect 3646 7588 3650 7644
rect 3650 7588 3706 7644
rect 3706 7588 3710 7644
rect 3646 7584 3710 7588
rect 3726 7644 3790 7648
rect 3726 7588 3730 7644
rect 3730 7588 3786 7644
rect 3786 7588 3790 7644
rect 3726 7584 3790 7588
rect 3806 7644 3870 7648
rect 3806 7588 3810 7644
rect 3810 7588 3866 7644
rect 3866 7588 3870 7644
rect 3806 7584 3870 7588
rect 3886 7644 3950 7648
rect 3886 7588 3890 7644
rect 3890 7588 3946 7644
rect 3946 7588 3950 7644
rect 3886 7584 3950 7588
rect 5002 7644 5066 7648
rect 5002 7588 5006 7644
rect 5006 7588 5062 7644
rect 5062 7588 5066 7644
rect 5002 7584 5066 7588
rect 5082 7644 5146 7648
rect 5082 7588 5086 7644
rect 5086 7588 5142 7644
rect 5142 7588 5146 7644
rect 5082 7584 5146 7588
rect 5162 7644 5226 7648
rect 5162 7588 5166 7644
rect 5166 7588 5222 7644
rect 5222 7588 5226 7644
rect 5162 7584 5226 7588
rect 5242 7644 5306 7648
rect 5242 7588 5246 7644
rect 5246 7588 5302 7644
rect 5302 7588 5306 7644
rect 5242 7584 5306 7588
rect 6358 7644 6422 7648
rect 6358 7588 6362 7644
rect 6362 7588 6418 7644
rect 6418 7588 6422 7644
rect 6358 7584 6422 7588
rect 6438 7644 6502 7648
rect 6438 7588 6442 7644
rect 6442 7588 6498 7644
rect 6498 7588 6502 7644
rect 6438 7584 6502 7588
rect 6518 7644 6582 7648
rect 6518 7588 6522 7644
rect 6522 7588 6578 7644
rect 6578 7588 6582 7644
rect 6518 7584 6582 7588
rect 6598 7644 6662 7648
rect 6598 7588 6602 7644
rect 6602 7588 6658 7644
rect 6658 7588 6662 7644
rect 6598 7584 6662 7588
rect 1630 7100 1694 7104
rect 1630 7044 1634 7100
rect 1634 7044 1690 7100
rect 1690 7044 1694 7100
rect 1630 7040 1694 7044
rect 1710 7100 1774 7104
rect 1710 7044 1714 7100
rect 1714 7044 1770 7100
rect 1770 7044 1774 7100
rect 1710 7040 1774 7044
rect 1790 7100 1854 7104
rect 1790 7044 1794 7100
rect 1794 7044 1850 7100
rect 1850 7044 1854 7100
rect 1790 7040 1854 7044
rect 1870 7100 1934 7104
rect 1870 7044 1874 7100
rect 1874 7044 1930 7100
rect 1930 7044 1934 7100
rect 1870 7040 1934 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 3146 7100 3210 7104
rect 3146 7044 3150 7100
rect 3150 7044 3206 7100
rect 3206 7044 3210 7100
rect 3146 7040 3210 7044
rect 3226 7100 3290 7104
rect 3226 7044 3230 7100
rect 3230 7044 3286 7100
rect 3286 7044 3290 7100
rect 3226 7040 3290 7044
rect 4342 7100 4406 7104
rect 4342 7044 4346 7100
rect 4346 7044 4402 7100
rect 4402 7044 4406 7100
rect 4342 7040 4406 7044
rect 4422 7100 4486 7104
rect 4422 7044 4426 7100
rect 4426 7044 4482 7100
rect 4482 7044 4486 7100
rect 4422 7040 4486 7044
rect 4502 7100 4566 7104
rect 4502 7044 4506 7100
rect 4506 7044 4562 7100
rect 4562 7044 4566 7100
rect 4502 7040 4566 7044
rect 4582 7100 4646 7104
rect 4582 7044 4586 7100
rect 4586 7044 4642 7100
rect 4642 7044 4646 7100
rect 4582 7040 4646 7044
rect 5698 7100 5762 7104
rect 5698 7044 5702 7100
rect 5702 7044 5758 7100
rect 5758 7044 5762 7100
rect 5698 7040 5762 7044
rect 5778 7100 5842 7104
rect 5778 7044 5782 7100
rect 5782 7044 5838 7100
rect 5838 7044 5842 7100
rect 5778 7040 5842 7044
rect 5858 7100 5922 7104
rect 5858 7044 5862 7100
rect 5862 7044 5918 7100
rect 5918 7044 5922 7100
rect 5858 7040 5922 7044
rect 5938 7100 6002 7104
rect 5938 7044 5942 7100
rect 5942 7044 5998 7100
rect 5998 7044 6002 7100
rect 5938 7040 6002 7044
rect 2290 6556 2354 6560
rect 2290 6500 2294 6556
rect 2294 6500 2350 6556
rect 2350 6500 2354 6556
rect 2290 6496 2354 6500
rect 2370 6556 2434 6560
rect 2370 6500 2374 6556
rect 2374 6500 2430 6556
rect 2430 6500 2434 6556
rect 2370 6496 2434 6500
rect 2450 6556 2514 6560
rect 2450 6500 2454 6556
rect 2454 6500 2510 6556
rect 2510 6500 2514 6556
rect 2450 6496 2514 6500
rect 2530 6556 2594 6560
rect 2530 6500 2534 6556
rect 2534 6500 2590 6556
rect 2590 6500 2594 6556
rect 2530 6496 2594 6500
rect 3646 6556 3710 6560
rect 3646 6500 3650 6556
rect 3650 6500 3706 6556
rect 3706 6500 3710 6556
rect 3646 6496 3710 6500
rect 3726 6556 3790 6560
rect 3726 6500 3730 6556
rect 3730 6500 3786 6556
rect 3786 6500 3790 6556
rect 3726 6496 3790 6500
rect 3806 6556 3870 6560
rect 3806 6500 3810 6556
rect 3810 6500 3866 6556
rect 3866 6500 3870 6556
rect 3806 6496 3870 6500
rect 3886 6556 3950 6560
rect 3886 6500 3890 6556
rect 3890 6500 3946 6556
rect 3946 6500 3950 6556
rect 3886 6496 3950 6500
rect 5002 6556 5066 6560
rect 5002 6500 5006 6556
rect 5006 6500 5062 6556
rect 5062 6500 5066 6556
rect 5002 6496 5066 6500
rect 5082 6556 5146 6560
rect 5082 6500 5086 6556
rect 5086 6500 5142 6556
rect 5142 6500 5146 6556
rect 5082 6496 5146 6500
rect 5162 6556 5226 6560
rect 5162 6500 5166 6556
rect 5166 6500 5222 6556
rect 5222 6500 5226 6556
rect 5162 6496 5226 6500
rect 5242 6556 5306 6560
rect 5242 6500 5246 6556
rect 5246 6500 5302 6556
rect 5302 6500 5306 6556
rect 5242 6496 5306 6500
rect 6358 6556 6422 6560
rect 6358 6500 6362 6556
rect 6362 6500 6418 6556
rect 6418 6500 6422 6556
rect 6358 6496 6422 6500
rect 6438 6556 6502 6560
rect 6438 6500 6442 6556
rect 6442 6500 6498 6556
rect 6498 6500 6502 6556
rect 6438 6496 6502 6500
rect 6518 6556 6582 6560
rect 6518 6500 6522 6556
rect 6522 6500 6578 6556
rect 6578 6500 6582 6556
rect 6518 6496 6582 6500
rect 6598 6556 6662 6560
rect 6598 6500 6602 6556
rect 6602 6500 6658 6556
rect 6658 6500 6662 6556
rect 6598 6496 6662 6500
rect 1630 6012 1694 6016
rect 1630 5956 1634 6012
rect 1634 5956 1690 6012
rect 1690 5956 1694 6012
rect 1630 5952 1694 5956
rect 1710 6012 1774 6016
rect 1710 5956 1714 6012
rect 1714 5956 1770 6012
rect 1770 5956 1774 6012
rect 1710 5952 1774 5956
rect 1790 6012 1854 6016
rect 1790 5956 1794 6012
rect 1794 5956 1850 6012
rect 1850 5956 1854 6012
rect 1790 5952 1854 5956
rect 1870 6012 1934 6016
rect 1870 5956 1874 6012
rect 1874 5956 1930 6012
rect 1930 5956 1934 6012
rect 1870 5952 1934 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 3146 6012 3210 6016
rect 3146 5956 3150 6012
rect 3150 5956 3206 6012
rect 3206 5956 3210 6012
rect 3146 5952 3210 5956
rect 3226 6012 3290 6016
rect 3226 5956 3230 6012
rect 3230 5956 3286 6012
rect 3286 5956 3290 6012
rect 3226 5952 3290 5956
rect 4342 6012 4406 6016
rect 4342 5956 4346 6012
rect 4346 5956 4402 6012
rect 4402 5956 4406 6012
rect 4342 5952 4406 5956
rect 4422 6012 4486 6016
rect 4422 5956 4426 6012
rect 4426 5956 4482 6012
rect 4482 5956 4486 6012
rect 4422 5952 4486 5956
rect 4502 6012 4566 6016
rect 4502 5956 4506 6012
rect 4506 5956 4562 6012
rect 4562 5956 4566 6012
rect 4502 5952 4566 5956
rect 4582 6012 4646 6016
rect 4582 5956 4586 6012
rect 4586 5956 4642 6012
rect 4642 5956 4646 6012
rect 4582 5952 4646 5956
rect 5698 6012 5762 6016
rect 5698 5956 5702 6012
rect 5702 5956 5758 6012
rect 5758 5956 5762 6012
rect 5698 5952 5762 5956
rect 5778 6012 5842 6016
rect 5778 5956 5782 6012
rect 5782 5956 5838 6012
rect 5838 5956 5842 6012
rect 5778 5952 5842 5956
rect 5858 6012 5922 6016
rect 5858 5956 5862 6012
rect 5862 5956 5918 6012
rect 5918 5956 5922 6012
rect 5858 5952 5922 5956
rect 5938 6012 6002 6016
rect 5938 5956 5942 6012
rect 5942 5956 5998 6012
rect 5998 5956 6002 6012
rect 5938 5952 6002 5956
rect 2290 5468 2354 5472
rect 2290 5412 2294 5468
rect 2294 5412 2350 5468
rect 2350 5412 2354 5468
rect 2290 5408 2354 5412
rect 2370 5468 2434 5472
rect 2370 5412 2374 5468
rect 2374 5412 2430 5468
rect 2430 5412 2434 5468
rect 2370 5408 2434 5412
rect 2450 5468 2514 5472
rect 2450 5412 2454 5468
rect 2454 5412 2510 5468
rect 2510 5412 2514 5468
rect 2450 5408 2514 5412
rect 2530 5468 2594 5472
rect 2530 5412 2534 5468
rect 2534 5412 2590 5468
rect 2590 5412 2594 5468
rect 2530 5408 2594 5412
rect 3646 5468 3710 5472
rect 3646 5412 3650 5468
rect 3650 5412 3706 5468
rect 3706 5412 3710 5468
rect 3646 5408 3710 5412
rect 3726 5468 3790 5472
rect 3726 5412 3730 5468
rect 3730 5412 3786 5468
rect 3786 5412 3790 5468
rect 3726 5408 3790 5412
rect 3806 5468 3870 5472
rect 3806 5412 3810 5468
rect 3810 5412 3866 5468
rect 3866 5412 3870 5468
rect 3806 5408 3870 5412
rect 3886 5468 3950 5472
rect 3886 5412 3890 5468
rect 3890 5412 3946 5468
rect 3946 5412 3950 5468
rect 3886 5408 3950 5412
rect 5002 5468 5066 5472
rect 5002 5412 5006 5468
rect 5006 5412 5062 5468
rect 5062 5412 5066 5468
rect 5002 5408 5066 5412
rect 5082 5468 5146 5472
rect 5082 5412 5086 5468
rect 5086 5412 5142 5468
rect 5142 5412 5146 5468
rect 5082 5408 5146 5412
rect 5162 5468 5226 5472
rect 5162 5412 5166 5468
rect 5166 5412 5222 5468
rect 5222 5412 5226 5468
rect 5162 5408 5226 5412
rect 5242 5468 5306 5472
rect 5242 5412 5246 5468
rect 5246 5412 5302 5468
rect 5302 5412 5306 5468
rect 5242 5408 5306 5412
rect 6358 5468 6422 5472
rect 6358 5412 6362 5468
rect 6362 5412 6418 5468
rect 6418 5412 6422 5468
rect 6358 5408 6422 5412
rect 6438 5468 6502 5472
rect 6438 5412 6442 5468
rect 6442 5412 6498 5468
rect 6498 5412 6502 5468
rect 6438 5408 6502 5412
rect 6518 5468 6582 5472
rect 6518 5412 6522 5468
rect 6522 5412 6578 5468
rect 6578 5412 6582 5468
rect 6518 5408 6582 5412
rect 6598 5468 6662 5472
rect 6598 5412 6602 5468
rect 6602 5412 6658 5468
rect 6658 5412 6662 5468
rect 6598 5408 6662 5412
rect 1630 4924 1694 4928
rect 1630 4868 1634 4924
rect 1634 4868 1690 4924
rect 1690 4868 1694 4924
rect 1630 4864 1694 4868
rect 1710 4924 1774 4928
rect 1710 4868 1714 4924
rect 1714 4868 1770 4924
rect 1770 4868 1774 4924
rect 1710 4864 1774 4868
rect 1790 4924 1854 4928
rect 1790 4868 1794 4924
rect 1794 4868 1850 4924
rect 1850 4868 1854 4924
rect 1790 4864 1854 4868
rect 1870 4924 1934 4928
rect 1870 4868 1874 4924
rect 1874 4868 1930 4924
rect 1930 4868 1934 4924
rect 1870 4864 1934 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 3146 4924 3210 4928
rect 3146 4868 3150 4924
rect 3150 4868 3206 4924
rect 3206 4868 3210 4924
rect 3146 4864 3210 4868
rect 3226 4924 3290 4928
rect 3226 4868 3230 4924
rect 3230 4868 3286 4924
rect 3286 4868 3290 4924
rect 3226 4864 3290 4868
rect 4342 4924 4406 4928
rect 4342 4868 4346 4924
rect 4346 4868 4402 4924
rect 4402 4868 4406 4924
rect 4342 4864 4406 4868
rect 4422 4924 4486 4928
rect 4422 4868 4426 4924
rect 4426 4868 4482 4924
rect 4482 4868 4486 4924
rect 4422 4864 4486 4868
rect 4502 4924 4566 4928
rect 4502 4868 4506 4924
rect 4506 4868 4562 4924
rect 4562 4868 4566 4924
rect 4502 4864 4566 4868
rect 4582 4924 4646 4928
rect 4582 4868 4586 4924
rect 4586 4868 4642 4924
rect 4642 4868 4646 4924
rect 4582 4864 4646 4868
rect 5698 4924 5762 4928
rect 5698 4868 5702 4924
rect 5702 4868 5758 4924
rect 5758 4868 5762 4924
rect 5698 4864 5762 4868
rect 5778 4924 5842 4928
rect 5778 4868 5782 4924
rect 5782 4868 5838 4924
rect 5838 4868 5842 4924
rect 5778 4864 5842 4868
rect 5858 4924 5922 4928
rect 5858 4868 5862 4924
rect 5862 4868 5918 4924
rect 5918 4868 5922 4924
rect 5858 4864 5922 4868
rect 5938 4924 6002 4928
rect 5938 4868 5942 4924
rect 5942 4868 5998 4924
rect 5998 4868 6002 4924
rect 5938 4864 6002 4868
rect 2290 4380 2354 4384
rect 2290 4324 2294 4380
rect 2294 4324 2350 4380
rect 2350 4324 2354 4380
rect 2290 4320 2354 4324
rect 2370 4380 2434 4384
rect 2370 4324 2374 4380
rect 2374 4324 2430 4380
rect 2430 4324 2434 4380
rect 2370 4320 2434 4324
rect 2450 4380 2514 4384
rect 2450 4324 2454 4380
rect 2454 4324 2510 4380
rect 2510 4324 2514 4380
rect 2450 4320 2514 4324
rect 2530 4380 2594 4384
rect 2530 4324 2534 4380
rect 2534 4324 2590 4380
rect 2590 4324 2594 4380
rect 2530 4320 2594 4324
rect 3646 4380 3710 4384
rect 3646 4324 3650 4380
rect 3650 4324 3706 4380
rect 3706 4324 3710 4380
rect 3646 4320 3710 4324
rect 3726 4380 3790 4384
rect 3726 4324 3730 4380
rect 3730 4324 3786 4380
rect 3786 4324 3790 4380
rect 3726 4320 3790 4324
rect 3806 4380 3870 4384
rect 3806 4324 3810 4380
rect 3810 4324 3866 4380
rect 3866 4324 3870 4380
rect 3806 4320 3870 4324
rect 3886 4380 3950 4384
rect 3886 4324 3890 4380
rect 3890 4324 3946 4380
rect 3946 4324 3950 4380
rect 3886 4320 3950 4324
rect 5002 4380 5066 4384
rect 5002 4324 5006 4380
rect 5006 4324 5062 4380
rect 5062 4324 5066 4380
rect 5002 4320 5066 4324
rect 5082 4380 5146 4384
rect 5082 4324 5086 4380
rect 5086 4324 5142 4380
rect 5142 4324 5146 4380
rect 5082 4320 5146 4324
rect 5162 4380 5226 4384
rect 5162 4324 5166 4380
rect 5166 4324 5222 4380
rect 5222 4324 5226 4380
rect 5162 4320 5226 4324
rect 5242 4380 5306 4384
rect 5242 4324 5246 4380
rect 5246 4324 5302 4380
rect 5302 4324 5306 4380
rect 5242 4320 5306 4324
rect 6358 4380 6422 4384
rect 6358 4324 6362 4380
rect 6362 4324 6418 4380
rect 6418 4324 6422 4380
rect 6358 4320 6422 4324
rect 6438 4380 6502 4384
rect 6438 4324 6442 4380
rect 6442 4324 6498 4380
rect 6498 4324 6502 4380
rect 6438 4320 6502 4324
rect 6518 4380 6582 4384
rect 6518 4324 6522 4380
rect 6522 4324 6578 4380
rect 6578 4324 6582 4380
rect 6518 4320 6582 4324
rect 6598 4380 6662 4384
rect 6598 4324 6602 4380
rect 6602 4324 6658 4380
rect 6658 4324 6662 4380
rect 6598 4320 6662 4324
rect 1630 3836 1694 3840
rect 1630 3780 1634 3836
rect 1634 3780 1690 3836
rect 1690 3780 1694 3836
rect 1630 3776 1694 3780
rect 1710 3836 1774 3840
rect 1710 3780 1714 3836
rect 1714 3780 1770 3836
rect 1770 3780 1774 3836
rect 1710 3776 1774 3780
rect 1790 3836 1854 3840
rect 1790 3780 1794 3836
rect 1794 3780 1850 3836
rect 1850 3780 1854 3836
rect 1790 3776 1854 3780
rect 1870 3836 1934 3840
rect 1870 3780 1874 3836
rect 1874 3780 1930 3836
rect 1930 3780 1934 3836
rect 1870 3776 1934 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 3146 3836 3210 3840
rect 3146 3780 3150 3836
rect 3150 3780 3206 3836
rect 3206 3780 3210 3836
rect 3146 3776 3210 3780
rect 3226 3836 3290 3840
rect 3226 3780 3230 3836
rect 3230 3780 3286 3836
rect 3286 3780 3290 3836
rect 3226 3776 3290 3780
rect 4342 3836 4406 3840
rect 4342 3780 4346 3836
rect 4346 3780 4402 3836
rect 4402 3780 4406 3836
rect 4342 3776 4406 3780
rect 4422 3836 4486 3840
rect 4422 3780 4426 3836
rect 4426 3780 4482 3836
rect 4482 3780 4486 3836
rect 4422 3776 4486 3780
rect 4502 3836 4566 3840
rect 4502 3780 4506 3836
rect 4506 3780 4562 3836
rect 4562 3780 4566 3836
rect 4502 3776 4566 3780
rect 4582 3836 4646 3840
rect 4582 3780 4586 3836
rect 4586 3780 4642 3836
rect 4642 3780 4646 3836
rect 4582 3776 4646 3780
rect 5698 3836 5762 3840
rect 5698 3780 5702 3836
rect 5702 3780 5758 3836
rect 5758 3780 5762 3836
rect 5698 3776 5762 3780
rect 5778 3836 5842 3840
rect 5778 3780 5782 3836
rect 5782 3780 5838 3836
rect 5838 3780 5842 3836
rect 5778 3776 5842 3780
rect 5858 3836 5922 3840
rect 5858 3780 5862 3836
rect 5862 3780 5918 3836
rect 5918 3780 5922 3836
rect 5858 3776 5922 3780
rect 5938 3836 6002 3840
rect 5938 3780 5942 3836
rect 5942 3780 5998 3836
rect 5998 3780 6002 3836
rect 5938 3776 6002 3780
rect 2290 3292 2354 3296
rect 2290 3236 2294 3292
rect 2294 3236 2350 3292
rect 2350 3236 2354 3292
rect 2290 3232 2354 3236
rect 2370 3292 2434 3296
rect 2370 3236 2374 3292
rect 2374 3236 2430 3292
rect 2430 3236 2434 3292
rect 2370 3232 2434 3236
rect 2450 3292 2514 3296
rect 2450 3236 2454 3292
rect 2454 3236 2510 3292
rect 2510 3236 2514 3292
rect 2450 3232 2514 3236
rect 2530 3292 2594 3296
rect 2530 3236 2534 3292
rect 2534 3236 2590 3292
rect 2590 3236 2594 3292
rect 2530 3232 2594 3236
rect 3646 3292 3710 3296
rect 3646 3236 3650 3292
rect 3650 3236 3706 3292
rect 3706 3236 3710 3292
rect 3646 3232 3710 3236
rect 3726 3292 3790 3296
rect 3726 3236 3730 3292
rect 3730 3236 3786 3292
rect 3786 3236 3790 3292
rect 3726 3232 3790 3236
rect 3806 3292 3870 3296
rect 3806 3236 3810 3292
rect 3810 3236 3866 3292
rect 3866 3236 3870 3292
rect 3806 3232 3870 3236
rect 3886 3292 3950 3296
rect 3886 3236 3890 3292
rect 3890 3236 3946 3292
rect 3946 3236 3950 3292
rect 3886 3232 3950 3236
rect 5002 3292 5066 3296
rect 5002 3236 5006 3292
rect 5006 3236 5062 3292
rect 5062 3236 5066 3292
rect 5002 3232 5066 3236
rect 5082 3292 5146 3296
rect 5082 3236 5086 3292
rect 5086 3236 5142 3292
rect 5142 3236 5146 3292
rect 5082 3232 5146 3236
rect 5162 3292 5226 3296
rect 5162 3236 5166 3292
rect 5166 3236 5222 3292
rect 5222 3236 5226 3292
rect 5162 3232 5226 3236
rect 5242 3292 5306 3296
rect 5242 3236 5246 3292
rect 5246 3236 5302 3292
rect 5302 3236 5306 3292
rect 5242 3232 5306 3236
rect 6358 3292 6422 3296
rect 6358 3236 6362 3292
rect 6362 3236 6418 3292
rect 6418 3236 6422 3292
rect 6358 3232 6422 3236
rect 6438 3292 6502 3296
rect 6438 3236 6442 3292
rect 6442 3236 6498 3292
rect 6498 3236 6502 3292
rect 6438 3232 6502 3236
rect 6518 3292 6582 3296
rect 6518 3236 6522 3292
rect 6522 3236 6578 3292
rect 6578 3236 6582 3292
rect 6518 3232 6582 3236
rect 6598 3292 6662 3296
rect 6598 3236 6602 3292
rect 6602 3236 6658 3292
rect 6658 3236 6662 3292
rect 6598 3232 6662 3236
rect 1630 2748 1694 2752
rect 1630 2692 1634 2748
rect 1634 2692 1690 2748
rect 1690 2692 1694 2748
rect 1630 2688 1694 2692
rect 1710 2748 1774 2752
rect 1710 2692 1714 2748
rect 1714 2692 1770 2748
rect 1770 2692 1774 2748
rect 1710 2688 1774 2692
rect 1790 2748 1854 2752
rect 1790 2692 1794 2748
rect 1794 2692 1850 2748
rect 1850 2692 1854 2748
rect 1790 2688 1854 2692
rect 1870 2748 1934 2752
rect 1870 2692 1874 2748
rect 1874 2692 1930 2748
rect 1930 2692 1934 2748
rect 1870 2688 1934 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 3146 2748 3210 2752
rect 3146 2692 3150 2748
rect 3150 2692 3206 2748
rect 3206 2692 3210 2748
rect 3146 2688 3210 2692
rect 3226 2748 3290 2752
rect 3226 2692 3230 2748
rect 3230 2692 3286 2748
rect 3286 2692 3290 2748
rect 3226 2688 3290 2692
rect 4342 2748 4406 2752
rect 4342 2692 4346 2748
rect 4346 2692 4402 2748
rect 4402 2692 4406 2748
rect 4342 2688 4406 2692
rect 4422 2748 4486 2752
rect 4422 2692 4426 2748
rect 4426 2692 4482 2748
rect 4482 2692 4486 2748
rect 4422 2688 4486 2692
rect 4502 2748 4566 2752
rect 4502 2692 4506 2748
rect 4506 2692 4562 2748
rect 4562 2692 4566 2748
rect 4502 2688 4566 2692
rect 4582 2748 4646 2752
rect 4582 2692 4586 2748
rect 4586 2692 4642 2748
rect 4642 2692 4646 2748
rect 4582 2688 4646 2692
rect 5698 2748 5762 2752
rect 5698 2692 5702 2748
rect 5702 2692 5758 2748
rect 5758 2692 5762 2748
rect 5698 2688 5762 2692
rect 5778 2748 5842 2752
rect 5778 2692 5782 2748
rect 5782 2692 5838 2748
rect 5838 2692 5842 2748
rect 5778 2688 5842 2692
rect 5858 2748 5922 2752
rect 5858 2692 5862 2748
rect 5862 2692 5918 2748
rect 5918 2692 5922 2748
rect 5858 2688 5922 2692
rect 5938 2748 6002 2752
rect 5938 2692 5942 2748
rect 5942 2692 5998 2748
rect 5998 2692 6002 2748
rect 5938 2688 6002 2692
rect 2290 2204 2354 2208
rect 2290 2148 2294 2204
rect 2294 2148 2350 2204
rect 2350 2148 2354 2204
rect 2290 2144 2354 2148
rect 2370 2204 2434 2208
rect 2370 2148 2374 2204
rect 2374 2148 2430 2204
rect 2430 2148 2434 2204
rect 2370 2144 2434 2148
rect 2450 2204 2514 2208
rect 2450 2148 2454 2204
rect 2454 2148 2510 2204
rect 2510 2148 2514 2204
rect 2450 2144 2514 2148
rect 2530 2204 2594 2208
rect 2530 2148 2534 2204
rect 2534 2148 2590 2204
rect 2590 2148 2594 2204
rect 2530 2144 2594 2148
rect 3646 2204 3710 2208
rect 3646 2148 3650 2204
rect 3650 2148 3706 2204
rect 3706 2148 3710 2204
rect 3646 2144 3710 2148
rect 3726 2204 3790 2208
rect 3726 2148 3730 2204
rect 3730 2148 3786 2204
rect 3786 2148 3790 2204
rect 3726 2144 3790 2148
rect 3806 2204 3870 2208
rect 3806 2148 3810 2204
rect 3810 2148 3866 2204
rect 3866 2148 3870 2204
rect 3806 2144 3870 2148
rect 3886 2204 3950 2208
rect 3886 2148 3890 2204
rect 3890 2148 3946 2204
rect 3946 2148 3950 2204
rect 3886 2144 3950 2148
rect 5002 2204 5066 2208
rect 5002 2148 5006 2204
rect 5006 2148 5062 2204
rect 5062 2148 5066 2204
rect 5002 2144 5066 2148
rect 5082 2204 5146 2208
rect 5082 2148 5086 2204
rect 5086 2148 5142 2204
rect 5142 2148 5146 2204
rect 5082 2144 5146 2148
rect 5162 2204 5226 2208
rect 5162 2148 5166 2204
rect 5166 2148 5222 2204
rect 5222 2148 5226 2204
rect 5162 2144 5226 2148
rect 5242 2204 5306 2208
rect 5242 2148 5246 2204
rect 5246 2148 5302 2204
rect 5302 2148 5306 2204
rect 5242 2144 5306 2148
rect 6358 2204 6422 2208
rect 6358 2148 6362 2204
rect 6362 2148 6418 2204
rect 6418 2148 6422 2204
rect 6358 2144 6422 2148
rect 6438 2204 6502 2208
rect 6438 2148 6442 2204
rect 6442 2148 6498 2204
rect 6498 2148 6502 2204
rect 6438 2144 6502 2148
rect 6518 2204 6582 2208
rect 6518 2148 6522 2204
rect 6522 2148 6578 2204
rect 6578 2148 6582 2204
rect 6518 2144 6582 2148
rect 6598 2204 6662 2208
rect 6598 2148 6602 2204
rect 6602 2148 6658 2204
rect 6658 2148 6662 2204
rect 6598 2144 6662 2148
<< metal4 >>
rect 1622 10368 1942 10384
rect 1622 10304 1630 10368
rect 1694 10304 1710 10368
rect 1774 10304 1790 10368
rect 1854 10304 1870 10368
rect 1934 10304 1942 10368
rect 1622 9434 1942 10304
rect 1622 9280 1664 9434
rect 1900 9280 1942 9434
rect 1622 9216 1630 9280
rect 1934 9216 1942 9280
rect 1622 9198 1664 9216
rect 1900 9198 1942 9216
rect 1622 8192 1942 9198
rect 1622 8128 1630 8192
rect 1694 8128 1710 8192
rect 1774 8128 1790 8192
rect 1854 8128 1870 8192
rect 1934 8128 1942 8192
rect 1622 7394 1942 8128
rect 1622 7158 1664 7394
rect 1900 7158 1942 7394
rect 1622 7104 1942 7158
rect 1622 7040 1630 7104
rect 1694 7040 1710 7104
rect 1774 7040 1790 7104
rect 1854 7040 1870 7104
rect 1934 7040 1942 7104
rect 1622 6016 1942 7040
rect 1622 5952 1630 6016
rect 1694 5952 1710 6016
rect 1774 5952 1790 6016
rect 1854 5952 1870 6016
rect 1934 5952 1942 6016
rect 1622 5354 1942 5952
rect 1622 5118 1664 5354
rect 1900 5118 1942 5354
rect 1622 4928 1942 5118
rect 1622 4864 1630 4928
rect 1694 4864 1710 4928
rect 1774 4864 1790 4928
rect 1854 4864 1870 4928
rect 1934 4864 1942 4928
rect 1622 3840 1942 4864
rect 1622 3776 1630 3840
rect 1694 3776 1710 3840
rect 1774 3776 1790 3840
rect 1854 3776 1870 3840
rect 1934 3776 1942 3840
rect 1622 3314 1942 3776
rect 1622 3078 1664 3314
rect 1900 3078 1942 3314
rect 1622 2752 1942 3078
rect 1622 2688 1630 2752
rect 1694 2688 1710 2752
rect 1774 2688 1790 2752
rect 1854 2688 1870 2752
rect 1934 2688 1942 2752
rect 1622 2128 1942 2688
rect 2282 10094 2602 10384
rect 2282 9858 2324 10094
rect 2560 9858 2602 10094
rect 2282 9824 2602 9858
rect 2282 9760 2290 9824
rect 2354 9760 2370 9824
rect 2434 9760 2450 9824
rect 2514 9760 2530 9824
rect 2594 9760 2602 9824
rect 2282 8736 2602 9760
rect 2282 8672 2290 8736
rect 2354 8672 2370 8736
rect 2434 8672 2450 8736
rect 2514 8672 2530 8736
rect 2594 8672 2602 8736
rect 2282 8054 2602 8672
rect 2282 7818 2324 8054
rect 2560 7818 2602 8054
rect 2282 7648 2602 7818
rect 2282 7584 2290 7648
rect 2354 7584 2370 7648
rect 2434 7584 2450 7648
rect 2514 7584 2530 7648
rect 2594 7584 2602 7648
rect 2282 6560 2602 7584
rect 2282 6496 2290 6560
rect 2354 6496 2370 6560
rect 2434 6496 2450 6560
rect 2514 6496 2530 6560
rect 2594 6496 2602 6560
rect 2282 6014 2602 6496
rect 2282 5778 2324 6014
rect 2560 5778 2602 6014
rect 2282 5472 2602 5778
rect 2282 5408 2290 5472
rect 2354 5408 2370 5472
rect 2434 5408 2450 5472
rect 2514 5408 2530 5472
rect 2594 5408 2602 5472
rect 2282 4384 2602 5408
rect 2282 4320 2290 4384
rect 2354 4320 2370 4384
rect 2434 4320 2450 4384
rect 2514 4320 2530 4384
rect 2594 4320 2602 4384
rect 2282 3974 2602 4320
rect 2282 3738 2324 3974
rect 2560 3738 2602 3974
rect 2282 3296 2602 3738
rect 2282 3232 2290 3296
rect 2354 3232 2370 3296
rect 2434 3232 2450 3296
rect 2514 3232 2530 3296
rect 2594 3232 2602 3296
rect 2282 2208 2602 3232
rect 2282 2144 2290 2208
rect 2354 2144 2370 2208
rect 2434 2144 2450 2208
rect 2514 2144 2530 2208
rect 2594 2144 2602 2208
rect 2282 2128 2602 2144
rect 2978 10368 3298 10384
rect 2978 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3146 10368
rect 3210 10304 3226 10368
rect 3290 10304 3298 10368
rect 2978 9434 3298 10304
rect 2978 9280 3020 9434
rect 3256 9280 3298 9434
rect 2978 9216 2986 9280
rect 3290 9216 3298 9280
rect 2978 9198 3020 9216
rect 3256 9198 3298 9216
rect 2978 8192 3298 9198
rect 2978 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3146 8192
rect 3210 8128 3226 8192
rect 3290 8128 3298 8192
rect 2978 7394 3298 8128
rect 2978 7158 3020 7394
rect 3256 7158 3298 7394
rect 2978 7104 3298 7158
rect 2978 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3146 7104
rect 3210 7040 3226 7104
rect 3290 7040 3298 7104
rect 2978 6016 3298 7040
rect 2978 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3146 6016
rect 3210 5952 3226 6016
rect 3290 5952 3298 6016
rect 2978 5354 3298 5952
rect 2978 5118 3020 5354
rect 3256 5118 3298 5354
rect 2978 4928 3298 5118
rect 2978 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3146 4928
rect 3210 4864 3226 4928
rect 3290 4864 3298 4928
rect 2978 3840 3298 4864
rect 2978 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3146 3840
rect 3210 3776 3226 3840
rect 3290 3776 3298 3840
rect 2978 3314 3298 3776
rect 2978 3078 3020 3314
rect 3256 3078 3298 3314
rect 2978 2752 3298 3078
rect 2978 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3146 2752
rect 3210 2688 3226 2752
rect 3290 2688 3298 2752
rect 2978 2128 3298 2688
rect 3638 10094 3958 10384
rect 3638 9858 3680 10094
rect 3916 9858 3958 10094
rect 3638 9824 3958 9858
rect 3638 9760 3646 9824
rect 3710 9760 3726 9824
rect 3790 9760 3806 9824
rect 3870 9760 3886 9824
rect 3950 9760 3958 9824
rect 3638 8736 3958 9760
rect 3638 8672 3646 8736
rect 3710 8672 3726 8736
rect 3790 8672 3806 8736
rect 3870 8672 3886 8736
rect 3950 8672 3958 8736
rect 3638 8054 3958 8672
rect 3638 7818 3680 8054
rect 3916 7818 3958 8054
rect 3638 7648 3958 7818
rect 3638 7584 3646 7648
rect 3710 7584 3726 7648
rect 3790 7584 3806 7648
rect 3870 7584 3886 7648
rect 3950 7584 3958 7648
rect 3638 6560 3958 7584
rect 3638 6496 3646 6560
rect 3710 6496 3726 6560
rect 3790 6496 3806 6560
rect 3870 6496 3886 6560
rect 3950 6496 3958 6560
rect 3638 6014 3958 6496
rect 3638 5778 3680 6014
rect 3916 5778 3958 6014
rect 3638 5472 3958 5778
rect 3638 5408 3646 5472
rect 3710 5408 3726 5472
rect 3790 5408 3806 5472
rect 3870 5408 3886 5472
rect 3950 5408 3958 5472
rect 3638 4384 3958 5408
rect 3638 4320 3646 4384
rect 3710 4320 3726 4384
rect 3790 4320 3806 4384
rect 3870 4320 3886 4384
rect 3950 4320 3958 4384
rect 3638 3974 3958 4320
rect 3638 3738 3680 3974
rect 3916 3738 3958 3974
rect 3638 3296 3958 3738
rect 3638 3232 3646 3296
rect 3710 3232 3726 3296
rect 3790 3232 3806 3296
rect 3870 3232 3886 3296
rect 3950 3232 3958 3296
rect 3638 2208 3958 3232
rect 3638 2144 3646 2208
rect 3710 2144 3726 2208
rect 3790 2144 3806 2208
rect 3870 2144 3886 2208
rect 3950 2144 3958 2208
rect 3638 2128 3958 2144
rect 4334 10368 4654 10384
rect 4334 10304 4342 10368
rect 4406 10304 4422 10368
rect 4486 10304 4502 10368
rect 4566 10304 4582 10368
rect 4646 10304 4654 10368
rect 4334 9434 4654 10304
rect 4334 9280 4376 9434
rect 4612 9280 4654 9434
rect 4334 9216 4342 9280
rect 4646 9216 4654 9280
rect 4334 9198 4376 9216
rect 4612 9198 4654 9216
rect 4334 8192 4654 9198
rect 4334 8128 4342 8192
rect 4406 8128 4422 8192
rect 4486 8128 4502 8192
rect 4566 8128 4582 8192
rect 4646 8128 4654 8192
rect 4334 7394 4654 8128
rect 4334 7158 4376 7394
rect 4612 7158 4654 7394
rect 4334 7104 4654 7158
rect 4334 7040 4342 7104
rect 4406 7040 4422 7104
rect 4486 7040 4502 7104
rect 4566 7040 4582 7104
rect 4646 7040 4654 7104
rect 4334 6016 4654 7040
rect 4334 5952 4342 6016
rect 4406 5952 4422 6016
rect 4486 5952 4502 6016
rect 4566 5952 4582 6016
rect 4646 5952 4654 6016
rect 4334 5354 4654 5952
rect 4334 5118 4376 5354
rect 4612 5118 4654 5354
rect 4334 4928 4654 5118
rect 4334 4864 4342 4928
rect 4406 4864 4422 4928
rect 4486 4864 4502 4928
rect 4566 4864 4582 4928
rect 4646 4864 4654 4928
rect 4334 3840 4654 4864
rect 4334 3776 4342 3840
rect 4406 3776 4422 3840
rect 4486 3776 4502 3840
rect 4566 3776 4582 3840
rect 4646 3776 4654 3840
rect 4334 3314 4654 3776
rect 4334 3078 4376 3314
rect 4612 3078 4654 3314
rect 4334 2752 4654 3078
rect 4334 2688 4342 2752
rect 4406 2688 4422 2752
rect 4486 2688 4502 2752
rect 4566 2688 4582 2752
rect 4646 2688 4654 2752
rect 4334 2128 4654 2688
rect 4994 10094 5314 10384
rect 4994 9858 5036 10094
rect 5272 9858 5314 10094
rect 4994 9824 5314 9858
rect 4994 9760 5002 9824
rect 5066 9760 5082 9824
rect 5146 9760 5162 9824
rect 5226 9760 5242 9824
rect 5306 9760 5314 9824
rect 4994 8736 5314 9760
rect 4994 8672 5002 8736
rect 5066 8672 5082 8736
rect 5146 8672 5162 8736
rect 5226 8672 5242 8736
rect 5306 8672 5314 8736
rect 4994 8054 5314 8672
rect 4994 7818 5036 8054
rect 5272 7818 5314 8054
rect 4994 7648 5314 7818
rect 4994 7584 5002 7648
rect 5066 7584 5082 7648
rect 5146 7584 5162 7648
rect 5226 7584 5242 7648
rect 5306 7584 5314 7648
rect 4994 6560 5314 7584
rect 4994 6496 5002 6560
rect 5066 6496 5082 6560
rect 5146 6496 5162 6560
rect 5226 6496 5242 6560
rect 5306 6496 5314 6560
rect 4994 6014 5314 6496
rect 4994 5778 5036 6014
rect 5272 5778 5314 6014
rect 4994 5472 5314 5778
rect 4994 5408 5002 5472
rect 5066 5408 5082 5472
rect 5146 5408 5162 5472
rect 5226 5408 5242 5472
rect 5306 5408 5314 5472
rect 4994 4384 5314 5408
rect 4994 4320 5002 4384
rect 5066 4320 5082 4384
rect 5146 4320 5162 4384
rect 5226 4320 5242 4384
rect 5306 4320 5314 4384
rect 4994 3974 5314 4320
rect 4994 3738 5036 3974
rect 5272 3738 5314 3974
rect 4994 3296 5314 3738
rect 4994 3232 5002 3296
rect 5066 3232 5082 3296
rect 5146 3232 5162 3296
rect 5226 3232 5242 3296
rect 5306 3232 5314 3296
rect 4994 2208 5314 3232
rect 4994 2144 5002 2208
rect 5066 2144 5082 2208
rect 5146 2144 5162 2208
rect 5226 2144 5242 2208
rect 5306 2144 5314 2208
rect 4994 2128 5314 2144
rect 5690 10368 6010 10384
rect 5690 10304 5698 10368
rect 5762 10304 5778 10368
rect 5842 10304 5858 10368
rect 5922 10304 5938 10368
rect 6002 10304 6010 10368
rect 5690 9434 6010 10304
rect 5690 9280 5732 9434
rect 5968 9280 6010 9434
rect 5690 9216 5698 9280
rect 6002 9216 6010 9280
rect 5690 9198 5732 9216
rect 5968 9198 6010 9216
rect 5690 8192 6010 9198
rect 5690 8128 5698 8192
rect 5762 8128 5778 8192
rect 5842 8128 5858 8192
rect 5922 8128 5938 8192
rect 6002 8128 6010 8192
rect 5690 7394 6010 8128
rect 5690 7158 5732 7394
rect 5968 7158 6010 7394
rect 5690 7104 6010 7158
rect 5690 7040 5698 7104
rect 5762 7040 5778 7104
rect 5842 7040 5858 7104
rect 5922 7040 5938 7104
rect 6002 7040 6010 7104
rect 5690 6016 6010 7040
rect 5690 5952 5698 6016
rect 5762 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5938 6016
rect 6002 5952 6010 6016
rect 5690 5354 6010 5952
rect 5690 5118 5732 5354
rect 5968 5118 6010 5354
rect 5690 4928 6010 5118
rect 5690 4864 5698 4928
rect 5762 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5938 4928
rect 6002 4864 6010 4928
rect 5690 3840 6010 4864
rect 5690 3776 5698 3840
rect 5762 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5938 3840
rect 6002 3776 6010 3840
rect 5690 3314 6010 3776
rect 5690 3078 5732 3314
rect 5968 3078 6010 3314
rect 5690 2752 6010 3078
rect 5690 2688 5698 2752
rect 5762 2688 5778 2752
rect 5842 2688 5858 2752
rect 5922 2688 5938 2752
rect 6002 2688 6010 2752
rect 5690 2128 6010 2688
rect 6350 10094 6670 10384
rect 6350 9858 6392 10094
rect 6628 9858 6670 10094
rect 6350 9824 6670 9858
rect 6350 9760 6358 9824
rect 6422 9760 6438 9824
rect 6502 9760 6518 9824
rect 6582 9760 6598 9824
rect 6662 9760 6670 9824
rect 6350 8736 6670 9760
rect 6350 8672 6358 8736
rect 6422 8672 6438 8736
rect 6502 8672 6518 8736
rect 6582 8672 6598 8736
rect 6662 8672 6670 8736
rect 6350 8054 6670 8672
rect 6350 7818 6392 8054
rect 6628 7818 6670 8054
rect 6350 7648 6670 7818
rect 6350 7584 6358 7648
rect 6422 7584 6438 7648
rect 6502 7584 6518 7648
rect 6582 7584 6598 7648
rect 6662 7584 6670 7648
rect 6350 6560 6670 7584
rect 6350 6496 6358 6560
rect 6422 6496 6438 6560
rect 6502 6496 6518 6560
rect 6582 6496 6598 6560
rect 6662 6496 6670 6560
rect 6350 6014 6670 6496
rect 6350 5778 6392 6014
rect 6628 5778 6670 6014
rect 6350 5472 6670 5778
rect 6350 5408 6358 5472
rect 6422 5408 6438 5472
rect 6502 5408 6518 5472
rect 6582 5408 6598 5472
rect 6662 5408 6670 5472
rect 6350 4384 6670 5408
rect 6350 4320 6358 4384
rect 6422 4320 6438 4384
rect 6502 4320 6518 4384
rect 6582 4320 6598 4384
rect 6662 4320 6670 4384
rect 6350 3974 6670 4320
rect 6350 3738 6392 3974
rect 6628 3738 6670 3974
rect 6350 3296 6670 3738
rect 6350 3232 6358 3296
rect 6422 3232 6438 3296
rect 6502 3232 6518 3296
rect 6582 3232 6598 3296
rect 6662 3232 6670 3296
rect 6350 2208 6670 3232
rect 6350 2144 6358 2208
rect 6422 2144 6438 2208
rect 6502 2144 6518 2208
rect 6582 2144 6598 2208
rect 6662 2144 6670 2208
rect 6350 2128 6670 2144
<< via4 >>
rect 1664 9280 1900 9434
rect 1664 9216 1694 9280
rect 1694 9216 1710 9280
rect 1710 9216 1774 9280
rect 1774 9216 1790 9280
rect 1790 9216 1854 9280
rect 1854 9216 1870 9280
rect 1870 9216 1900 9280
rect 1664 9198 1900 9216
rect 1664 7158 1900 7394
rect 1664 5118 1900 5354
rect 1664 3078 1900 3314
rect 2324 9858 2560 10094
rect 2324 7818 2560 8054
rect 2324 5778 2560 6014
rect 2324 3738 2560 3974
rect 3020 9280 3256 9434
rect 3020 9216 3050 9280
rect 3050 9216 3066 9280
rect 3066 9216 3130 9280
rect 3130 9216 3146 9280
rect 3146 9216 3210 9280
rect 3210 9216 3226 9280
rect 3226 9216 3256 9280
rect 3020 9198 3256 9216
rect 3020 7158 3256 7394
rect 3020 5118 3256 5354
rect 3020 3078 3256 3314
rect 3680 9858 3916 10094
rect 3680 7818 3916 8054
rect 3680 5778 3916 6014
rect 3680 3738 3916 3974
rect 4376 9280 4612 9434
rect 4376 9216 4406 9280
rect 4406 9216 4422 9280
rect 4422 9216 4486 9280
rect 4486 9216 4502 9280
rect 4502 9216 4566 9280
rect 4566 9216 4582 9280
rect 4582 9216 4612 9280
rect 4376 9198 4612 9216
rect 4376 7158 4612 7394
rect 4376 5118 4612 5354
rect 4376 3078 4612 3314
rect 5036 9858 5272 10094
rect 5036 7818 5272 8054
rect 5036 5778 5272 6014
rect 5036 3738 5272 3974
rect 5732 9280 5968 9434
rect 5732 9216 5762 9280
rect 5762 9216 5778 9280
rect 5778 9216 5842 9280
rect 5842 9216 5858 9280
rect 5858 9216 5922 9280
rect 5922 9216 5938 9280
rect 5938 9216 5968 9280
rect 5732 9198 5968 9216
rect 5732 7158 5968 7394
rect 5732 5118 5968 5354
rect 5732 3078 5968 3314
rect 6392 9858 6628 10094
rect 6392 7818 6628 8054
rect 6392 5778 6628 6014
rect 6392 3738 6628 3974
<< metal5 >>
rect 1056 10094 6670 10136
rect 1056 9858 2324 10094
rect 2560 9858 3680 10094
rect 3916 9858 5036 10094
rect 5272 9858 6392 10094
rect 6628 9858 6670 10094
rect 1056 9816 6670 9858
rect 1056 9434 6580 9476
rect 1056 9198 1664 9434
rect 1900 9198 3020 9434
rect 3256 9198 4376 9434
rect 4612 9198 5732 9434
rect 5968 9198 6580 9434
rect 1056 9156 6580 9198
rect 1056 8054 6670 8096
rect 1056 7818 2324 8054
rect 2560 7818 3680 8054
rect 3916 7818 5036 8054
rect 5272 7818 6392 8054
rect 6628 7818 6670 8054
rect 1056 7776 6670 7818
rect 1056 7394 6580 7436
rect 1056 7158 1664 7394
rect 1900 7158 3020 7394
rect 3256 7158 4376 7394
rect 4612 7158 5732 7394
rect 5968 7158 6580 7394
rect 1056 7116 6580 7158
rect 1056 6014 6670 6056
rect 1056 5778 2324 6014
rect 2560 5778 3680 6014
rect 3916 5778 5036 6014
rect 5272 5778 6392 6014
rect 6628 5778 6670 6014
rect 1056 5736 6670 5778
rect 1056 5354 6580 5396
rect 1056 5118 1664 5354
rect 1900 5118 3020 5354
rect 3256 5118 4376 5354
rect 4612 5118 5732 5354
rect 5968 5118 6580 5354
rect 1056 5076 6580 5118
rect 1056 3974 6670 4016
rect 1056 3738 2324 3974
rect 2560 3738 3680 3974
rect 3916 3738 5036 3974
rect 5272 3738 6392 3974
rect 6628 3738 6670 3974
rect 1056 3696 6670 3738
rect 1056 3314 6580 3356
rect 1056 3078 1664 3314
rect 1900 3078 3020 3314
rect 3256 3078 4376 3314
rect 4612 3078 5732 3314
rect 5968 3078 6580 3314
rect 1056 3036 6580 3078
use sky130_fd_sc_hd__buf_2  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1564 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _34_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1932 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _35_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1701704242
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 3496 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3772 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1701704242
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _40_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3312 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _42_
timestamp 1701704242
transform -1 0 4416 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _43_
timestamp 1701704242
transform -1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _44_
timestamp 1701704242
transform -1 0 6072 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _45_
timestamp 1701704242
transform 1 0 4324 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _46_
timestamp 1701704242
transform 1 0 5060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _47_
timestamp 1701704242
transform 1 0 4692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _48_
timestamp 1701704242
transform -1 0 6072 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _49_
timestamp 1701704242
transform 1 0 4416 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _50_
timestamp 1701704242
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _51_
timestamp 1701704242
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _52_
timestamp 1701704242
transform -1 0 4784 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _53_
timestamp 1701704242
transform 1 0 3220 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _54_
timestamp 1701704242
transform -1 0 2576 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _55_
timestamp 1701704242
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _56_
timestamp 1701704242
transform -1 0 3864 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _57_
timestamp 1701704242
transform 1 0 2576 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _58_
timestamp 1701704242
transform 1 0 4600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _59_
timestamp 1701704242
transform 1 0 3864 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _60_
timestamp 1701704242
transform 1 0 3220 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _61_
timestamp 1701704242
transform -1 0 4600 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _62_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _63_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _64_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1472 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _65_
timestamp 1701704242
transform -1 0 3404 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _66_
timestamp 1701704242
transform 1 0 4324 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _67_
timestamp 1701704242
transform 1 0 4324 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _68_
timestamp 1701704242
transform -1 0 3220 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _69_
timestamp 1701704242
transform -1 0 3404 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _70_
timestamp 1701704242
transform 1 0 4140 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _71_
timestamp 1701704242
transform 1 0 4416 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _72_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1701704242
transform 1 0 3772 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1701704242
transform -1 0 4416 0 -1 8704
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_45
timestamp 1701704242
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 2300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_42
timestamp 1701704242
transform 1 0 4968 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1701704242
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 1701704242
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_54
timestamp 1701704242
transform 1 0 6072 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1701704242
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_31
timestamp 1701704242
transform 1 0 3956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_25
timestamp 1701704242
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_55
timestamp 1701704242
transform 1 0 6164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1701704242
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_19
timestamp 1701704242
transform 1 0 2852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1701704242
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 1701704242
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1701704242
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1701704242
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_35
timestamp 1701704242
transform 1 0 4324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_45
timestamp 1701704242
transform 1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_49
timestamp 1701704242
transform 1 0 5612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_6
timestamp 1701704242
transform 1 0 1656 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_14
timestamp 1701704242
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_20
timestamp 1701704242
transform 1 0 2944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_45
timestamp 1701704242
transform 1 0 5244 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_51
timestamp 1701704242
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1701704242
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_40
timestamp 1701704242
transform 1 0 4784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_48
timestamp 1701704242
transform 1 0 5520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_30
timestamp 1701704242
transform 1 0 3864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_44
timestamp 1701704242
transform 1 0 5152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1701704242
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 1701704242
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_53
timestamp 1701704242
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_15
timestamp 1701704242
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1701704242
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_15
timestamp 1701704242
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_21
timestamp 1701704242
transform 1 0 3036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_36
timestamp 1701704242
transform 1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_9
timestamp 1701704242
transform 1 0 1932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_21
timestamp 1701704242
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_30
timestamp 1701704242
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_42
timestamp 1701704242
transform 1 0 4968 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_51
timestamp 1701704242
transform 1 0 5796 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_7
timestamp 1701704242
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1701704242
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_41
timestamp 1701704242
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_54
timestamp 1701704242
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1701704242
transform -1 0 5520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1701704242
transform -1 0 3404 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1701704242
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1701704242
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1701704242
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1701704242
transform 1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1701704242
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1701704242
transform 1 0 5704 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1701704242
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1701704242
transform 1 0 5704 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1701704242
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1701704242
transform 1 0 5152 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1701704242
transform 1 0 5520 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_15
timestamp 1701704242
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_16
timestamp 1701704242
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_17
timestamp 1701704242
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_18
timestamp 1701704242
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_19
timestamp 1701704242
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_20
timestamp 1701704242
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_21
timestamp 1701704242
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_22
timestamp 1701704242
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_23
timestamp 1701704242
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_24
timestamp 1701704242
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_25
timestamp 1701704242
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_26
timestamp 1701704242
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_27
timestamp 1701704242
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_28
timestamp 1701704242
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_29
timestamp 1701704242
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 6532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_31
timestamp 1701704242
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_32
timestamp 1701704242
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_33
timestamp 1701704242
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_34
timestamp 1701704242
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_35
timestamp 1701704242
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_36
timestamp 1701704242
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_37
timestamp 1701704242
transform 1 0 3680 0 1 9792
box -38 -48 130 592
<< labels >>
flabel metal4 s 2282 2128 2602 10384 0 FreeSans 1920 90 0 0 GND
port 0 nsew ground bidirectional
flabel metal4 s 3638 2128 3958 10384 0 FreeSans 1920 90 0 0 GND
port 0 nsew ground bidirectional
flabel metal4 s 4994 2128 5314 10384 0 FreeSans 1920 90 0 0 GND
port 0 nsew ground bidirectional
flabel metal4 s 6350 2128 6670 10384 0 FreeSans 1920 90 0 0 GND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3696 6670 4016 0 FreeSans 2560 0 0 0 GND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5736 6670 6056 0 FreeSans 2560 0 0 0 GND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7776 6670 8096 0 FreeSans 2560 0 0 0 GND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9816 6670 10136 0 FreeSans 2560 0 0 0 GND
port 0 nsew ground bidirectional
flabel metal4 s 1622 2128 1942 10384 0 FreeSans 1920 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 2978 2128 3298 10384 0 FreeSans 1920 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 4334 2128 4654 10384 0 FreeSans 1920 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 5690 2128 6010 10384 0 FreeSans 1920 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal5 s 1056 3036 6580 3356 0 FreeSans 2560 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal5 s 1056 5076 6580 5396 0 FreeSans 2560 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal5 s 1056 7116 6580 7436 0 FreeSans 2560 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal5 s 1056 9156 6580 9476 0 FreeSans 2560 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 6901 552 7701 672 0 FreeSans 480 0 0 0 data_out[0]
port 3 nsew signal tristate
flabel metal3 s 6901 1912 7701 2032 0 FreeSans 480 0 0 0 data_out[1]
port 4 nsew signal tristate
flabel metal3 s 6901 3272 7701 3392 0 FreeSans 480 0 0 0 data_out[2]
port 5 nsew signal tristate
flabel metal3 s 6901 4632 7701 4752 0 FreeSans 480 0 0 0 data_out[3]
port 6 nsew signal tristate
flabel metal3 s 6901 5992 7701 6112 0 FreeSans 480 0 0 0 data_out[4]
port 7 nsew signal tristate
flabel metal3 s 6901 7352 7701 7472 0 FreeSans 480 0 0 0 data_out[5]
port 8 nsew signal tristate
flabel metal3 s 6901 8712 7701 8832 0 FreeSans 480 0 0 0 data_out[6]
port 9 nsew signal tristate
flabel metal3 s 6901 10072 7701 10192 0 FreeSans 480 0 0 0 data_out[7]
port 10 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 enable
port 11 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 reset
port 12 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 scan_en
port 13 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 scan_in
port 14 nsew signal input
flabel metal3 s 6901 11432 7701 11552 0 FreeSans 480 0 0 0 scan_out
port 15 nsew signal tristate
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 shift
port 16 nsew signal input
rlabel via1 3887 9792 3887 9792 0 GND
rlabel metal1 3818 10336 3818 10336 0 VDD
rlabel metal1 1840 4046 1840 4046 0 _00_
rlabel metal1 3220 3434 3220 3434 0 _01_
rlabel metal1 4554 3162 4554 3162 0 _02_
rlabel metal1 4830 4658 4830 4658 0 _03_
rlabel metal1 3082 7310 3082 7310 0 _04_
rlabel metal2 2806 7378 2806 7378 0 _05_
rlabel metal1 4508 7514 4508 7514 0 _06_
rlabel metal1 5520 9010 5520 9010 0 _07_
rlabel metal1 5750 8976 5750 8976 0 _08_
rlabel metal1 3542 4148 3542 4148 0 _09_
rlabel metal1 2622 4607 2622 4607 0 _10_
rlabel metal1 4094 9010 4094 9010 0 _11_
rlabel metal1 3542 4046 3542 4046 0 _12_
rlabel metal1 3910 3162 3910 3162 0 _13_
rlabel metal1 5106 7378 5106 7378 0 _14_
rlabel metal1 3496 3162 3496 3162 0 _15_
rlabel metal1 4738 2890 4738 2890 0 _16_
rlabel metal1 4508 2958 4508 2958 0 _17_
rlabel metal1 5124 3026 5124 3026 0 _18_
rlabel metal1 4922 5134 4922 5134 0 _19_
rlabel metal1 4784 5202 4784 5202 0 _20_
rlabel metal1 5612 3706 5612 3706 0 _21_
rlabel metal1 3680 5882 3680 5882 0 _22_
rlabel metal1 3726 6970 3726 6970 0 _23_
rlabel metal1 4324 6970 4324 6970 0 _24_
rlabel metal1 2714 6834 2714 6834 0 _25_
rlabel via1 2990 6851 2990 6851 0 _26_
rlabel metal1 3082 6800 3082 6800 0 _27_
rlabel metal1 4462 7242 4462 7242 0 _28_
rlabel metal1 4186 7208 4186 7208 0 _29_
rlabel metal1 3864 6630 3864 6630 0 _30_
rlabel metal1 6210 9010 6210 9010 0 _31_
rlabel metal3 1740 1428 1740 1428 0 clk
rlabel metal1 4278 6086 4278 6086 0 clknet_0_clk
rlabel metal2 1518 3876 1518 3876 0 clknet_1_0__leaf_clk
rlabel metal2 3358 8092 3358 8092 0 clknet_1_1__leaf_clk
rlabel metal1 6164 2278 6164 2278 0 data_out[0]
rlabel metal2 5566 2125 5566 2125 0 data_out[1]
rlabel metal1 6440 3162 6440 3162 0 data_out[2]
rlabel metal1 6164 5542 6164 5542 0 data_out[3]
rlabel via2 6118 6069 6118 6069 0 data_out[4]
rlabel metal1 6164 6834 6164 6834 0 data_out[5]
rlabel metal1 6440 9350 6440 9350 0 data_out[6]
rlabel metal2 5382 10183 5382 10183 0 data_out[7]
rlabel metal3 820 10948 820 10948 0 enable
rlabel metal1 2576 9894 2576 9894 0 net1
rlabel metal1 2300 6766 2300 6766 0 net10
rlabel metal1 4232 6834 4232 6834 0 net11
rlabel metal2 3542 8500 3542 8500 0 net12
rlabel metal1 5934 8908 5934 8908 0 net13
rlabel metal2 5382 9826 5382 9826 0 net14
rlabel metal1 6164 7514 6164 7514 0 net15
rlabel metal1 4784 8398 4784 8398 0 net16
rlabel metal1 2530 4522 2530 4522 0 net17
rlabel metal2 1978 8602 1978 8602 0 net2
rlabel metal1 3358 6732 3358 6732 0 net3
rlabel metal1 2047 4590 2047 4590 0 net4
rlabel metal1 1702 5270 1702 5270 0 net5
rlabel metal1 4968 2346 4968 2346 0 net6
rlabel metal1 3082 2992 3082 2992 0 net7
rlabel metal1 5934 3060 5934 3060 0 net8
rlabel metal1 6164 4454 6164 4454 0 net9
rlabel metal3 820 9044 820 9044 0 reset
rlabel metal3 751 7140 751 7140 0 scan_en
rlabel metal3 1050 5236 1050 5236 0 scan_in
rlabel metal1 6164 10234 6164 10234 0 scan_out
rlabel metal3 820 3332 820 3332 0 shift
<< properties >>
string FIXED_BBOX 0 0 7701 12592
<< end >>
