magic
tech sky130A
magscale 1 2
timestamp 1698611618
<< error_p >>
rect -554 123 -496 129
rect -554 89 -542 123
rect -218 104 -158 142
rect -134 123 -76 129
rect -134 89 -122 123
rect 202 104 262 142
rect 286 123 344 129
rect 286 89 298 123
rect 622 104 682 142
rect 706 123 764 129
rect 706 89 718 123
rect -554 83 -496 89
rect -134 83 -76 89
rect 286 83 344 89
rect 706 83 764 89
rect -764 -89 -706 -83
rect -344 -89 -286 -83
rect 76 -89 134 -83
rect 496 -89 554 -83
rect -764 -123 -752 -89
rect -764 -129 -706 -123
rect -428 -142 -368 -104
rect -344 -123 -332 -89
rect -344 -129 -286 -123
rect -8 -142 52 -104
rect 76 -123 88 -89
rect 76 -129 134 -123
rect 412 -142 472 -104
rect 496 -123 508 -89
rect 496 -129 554 -123
<< nwell >>
rect -638 104 -412 142
rect -218 104 8 142
rect 202 104 428 142
rect 622 104 848 142
rect -848 -104 848 104
rect -848 -142 -622 -104
rect -428 -142 -202 -104
rect -8 -142 218 -104
rect 412 -142 638 -104
<< pmos >>
rect -750 -42 -720 42
rect -540 -42 -510 42
rect -330 -42 -300 42
rect -120 -42 -90 42
rect 90 -42 120 42
rect 300 -42 330 42
rect 510 -42 540 42
rect 720 -42 750 42
<< pdiff >>
rect -812 30 -750 42
rect -812 -30 -800 30
rect -766 -30 -750 30
rect -812 -42 -750 -30
rect -720 30 -658 42
rect -720 -30 -704 30
rect -670 -30 -658 30
rect -720 -42 -658 -30
rect -602 30 -540 42
rect -602 -30 -590 30
rect -556 -30 -540 30
rect -602 -42 -540 -30
rect -510 30 -448 42
rect -510 -30 -494 30
rect -460 -30 -448 30
rect -510 -42 -448 -30
rect -392 30 -330 42
rect -392 -30 -380 30
rect -346 -30 -330 30
rect -392 -42 -330 -30
rect -300 30 -238 42
rect -300 -30 -284 30
rect -250 -30 -238 30
rect -300 -42 -238 -30
rect -182 30 -120 42
rect -182 -30 -170 30
rect -136 -30 -120 30
rect -182 -42 -120 -30
rect -90 30 -28 42
rect -90 -30 -74 30
rect -40 -30 -28 30
rect -90 -42 -28 -30
rect 28 30 90 42
rect 28 -30 40 30
rect 74 -30 90 30
rect 28 -42 90 -30
rect 120 30 182 42
rect 120 -30 136 30
rect 170 -30 182 30
rect 120 -42 182 -30
rect 238 30 300 42
rect 238 -30 250 30
rect 284 -30 300 30
rect 238 -42 300 -30
rect 330 30 392 42
rect 330 -30 346 30
rect 380 -30 392 30
rect 330 -42 392 -30
rect 448 30 510 42
rect 448 -30 460 30
rect 494 -30 510 30
rect 448 -42 510 -30
rect 540 30 602 42
rect 540 -30 556 30
rect 590 -30 602 30
rect 540 -42 602 -30
rect 658 30 720 42
rect 658 -30 670 30
rect 704 -30 720 30
rect 658 -42 720 -30
rect 750 30 812 42
rect 750 -30 766 30
rect 800 -30 812 30
rect 750 -42 812 -30
<< pdiffc >>
rect -800 -30 -766 30
rect -704 -30 -670 30
rect -590 -30 -556 30
rect -494 -30 -460 30
rect -380 -30 -346 30
rect -284 -30 -250 30
rect -170 -30 -136 30
rect -74 -30 -40 30
rect 40 -30 74 30
rect 136 -30 170 30
rect 250 -30 284 30
rect 346 -30 380 30
rect 460 -30 494 30
rect 556 -30 590 30
rect 670 -30 704 30
rect 766 -30 800 30
<< poly >>
rect -558 123 -492 139
rect -558 89 -542 123
rect -508 89 -492 123
rect -558 73 -492 89
rect -138 123 -72 139
rect -138 89 -122 123
rect -88 89 -72 123
rect -138 73 -72 89
rect 282 123 348 139
rect 282 89 298 123
rect 332 89 348 123
rect 282 73 348 89
rect 702 123 768 139
rect 702 89 718 123
rect 752 89 768 123
rect 702 73 768 89
rect -750 42 -720 68
rect -540 42 -510 73
rect -330 42 -300 68
rect -120 42 -90 73
rect 90 42 120 68
rect 300 42 330 73
rect 510 42 540 68
rect 720 42 750 73
rect -750 -73 -720 -42
rect -540 -68 -510 -42
rect -330 -73 -300 -42
rect -120 -68 -90 -42
rect 90 -73 120 -42
rect 300 -68 330 -42
rect 510 -73 540 -42
rect 720 -68 750 -42
rect -768 -89 -702 -73
rect -768 -123 -752 -89
rect -718 -123 -702 -89
rect -768 -139 -702 -123
rect -348 -89 -282 -73
rect -348 -123 -332 -89
rect -298 -123 -282 -89
rect -348 -139 -282 -123
rect 72 -89 138 -73
rect 72 -123 88 -89
rect 122 -123 138 -89
rect 72 -139 138 -123
rect 492 -89 558 -73
rect 492 -123 508 -89
rect 542 -123 558 -89
rect 492 -139 558 -123
<< polycont >>
rect -542 89 -508 123
rect -122 89 -88 123
rect 298 89 332 123
rect 718 89 752 123
rect -752 -123 -718 -89
rect -332 -123 -298 -89
rect 88 -123 122 -89
rect 508 -123 542 -89
<< locali >>
rect -558 89 -542 123
rect -508 89 -492 123
rect -138 89 -122 123
rect -88 89 -72 123
rect 282 89 298 123
rect 332 89 348 123
rect 702 89 718 123
rect 752 89 768 123
rect -800 30 -766 46
rect -800 -46 -766 -30
rect -704 30 -670 46
rect -704 -46 -670 -30
rect -590 30 -556 46
rect -590 -46 -556 -30
rect -494 30 -460 46
rect -494 -46 -460 -30
rect -380 30 -346 46
rect -380 -46 -346 -30
rect -284 30 -250 46
rect -284 -46 -250 -30
rect -170 30 -136 46
rect -170 -46 -136 -30
rect -74 30 -40 46
rect -74 -46 -40 -30
rect 40 30 74 46
rect 40 -46 74 -30
rect 136 30 170 46
rect 136 -46 170 -30
rect 250 30 284 46
rect 250 -46 284 -30
rect 346 30 380 46
rect 346 -46 380 -30
rect 460 30 494 46
rect 460 -46 494 -30
rect 556 30 590 46
rect 556 -46 590 -30
rect 670 30 704 46
rect 670 -46 704 -30
rect 766 30 800 46
rect 766 -46 800 -30
rect -768 -123 -752 -89
rect -718 -123 -702 -89
rect -348 -123 -332 -89
rect -298 -123 -282 -89
rect 72 -123 88 -89
rect 122 -123 138 -89
rect 492 -123 508 -89
rect 542 -123 558 -89
<< viali >>
rect -542 89 -508 123
rect -122 89 -88 123
rect 298 89 332 123
rect 718 89 752 123
rect -800 -30 -766 30
rect -704 -30 -670 30
rect -590 -30 -556 30
rect -494 -30 -460 30
rect -380 -30 -346 30
rect -284 -30 -250 30
rect -170 -30 -136 30
rect -74 -30 -40 30
rect 40 -30 74 30
rect 136 -30 170 30
rect 250 -30 284 30
rect 346 -30 380 30
rect 460 -30 494 30
rect 556 -30 590 30
rect 670 -30 704 30
rect 766 -30 800 30
rect -752 -123 -718 -89
rect -332 -123 -298 -89
rect 88 -123 122 -89
rect 508 -123 542 -89
<< metal1 >>
rect -554 123 -496 129
rect -554 89 -542 123
rect -508 89 -496 123
rect -554 83 -496 89
rect -134 123 -76 129
rect -134 89 -122 123
rect -88 89 -76 123
rect -134 83 -76 89
rect 286 123 344 129
rect 286 89 298 123
rect 332 89 344 123
rect 286 83 344 89
rect 706 123 764 129
rect 706 89 718 123
rect 752 89 764 123
rect 706 83 764 89
rect -806 30 -760 42
rect -806 -30 -800 30
rect -766 -30 -760 30
rect -806 -42 -760 -30
rect -710 30 -664 42
rect -710 -30 -704 30
rect -670 -30 -664 30
rect -710 -42 -664 -30
rect -596 30 -550 42
rect -596 -30 -590 30
rect -556 -30 -550 30
rect -596 -42 -550 -30
rect -500 30 -454 42
rect -500 -30 -494 30
rect -460 -30 -454 30
rect -500 -42 -454 -30
rect -386 30 -340 42
rect -386 -30 -380 30
rect -346 -30 -340 30
rect -386 -42 -340 -30
rect -290 30 -244 42
rect -290 -30 -284 30
rect -250 -30 -244 30
rect -290 -42 -244 -30
rect -176 30 -130 42
rect -176 -30 -170 30
rect -136 -30 -130 30
rect -176 -42 -130 -30
rect -80 30 -34 42
rect -80 -30 -74 30
rect -40 -30 -34 30
rect -80 -42 -34 -30
rect 34 30 80 42
rect 34 -30 40 30
rect 74 -30 80 30
rect 34 -42 80 -30
rect 130 30 176 42
rect 130 -30 136 30
rect 170 -30 176 30
rect 130 -42 176 -30
rect 244 30 290 42
rect 244 -30 250 30
rect 284 -30 290 30
rect 244 -42 290 -30
rect 340 30 386 42
rect 340 -30 346 30
rect 380 -30 386 30
rect 340 -42 386 -30
rect 454 30 500 42
rect 454 -30 460 30
rect 494 -30 500 30
rect 454 -42 500 -30
rect 550 30 596 42
rect 550 -30 556 30
rect 590 -30 596 30
rect 550 -42 596 -30
rect 664 30 710 42
rect 664 -30 670 30
rect 704 -30 710 30
rect 664 -42 710 -30
rect 760 30 806 42
rect 760 -30 766 30
rect 800 -30 806 30
rect 760 -42 806 -30
rect -764 -89 -706 -83
rect -764 -123 -752 -89
rect -718 -123 -706 -89
rect -764 -129 -706 -123
rect -344 -89 -286 -83
rect -344 -123 -332 -89
rect -298 -123 -286 -89
rect -344 -129 -286 -123
rect 76 -89 134 -83
rect 76 -123 88 -89
rect 122 -123 134 -89
rect 76 -129 134 -123
rect 496 -89 554 -83
rect 496 -123 508 -89
rect 542 -123 554 -89
rect 496 -129 554 -123
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
