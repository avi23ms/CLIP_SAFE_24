magic
tech sky130A
magscale 1 2
timestamp 1697915631
<< pwell >>
rect -641 -252 641 252
<< nmos >>
rect -445 -42 -345 42
rect -287 -42 -187 42
rect -129 -42 -29 42
rect 29 -42 129 42
rect 187 -42 287 42
rect 345 -42 445 42
<< ndiff >>
rect -503 30 -445 42
rect -503 -30 -491 30
rect -457 -30 -445 30
rect -503 -42 -445 -30
rect -345 30 -287 42
rect -345 -30 -333 30
rect -299 -30 -287 30
rect -345 -42 -287 -30
rect -187 30 -129 42
rect -187 -30 -175 30
rect -141 -30 -129 30
rect -187 -42 -129 -30
rect -29 30 29 42
rect -29 -30 -17 30
rect 17 -30 29 30
rect -29 -42 29 -30
rect 129 30 187 42
rect 129 -30 141 30
rect 175 -30 187 30
rect 129 -42 187 -30
rect 287 30 345 42
rect 287 -30 299 30
rect 333 -30 345 30
rect 287 -42 345 -30
rect 445 30 503 42
rect 445 -30 457 30
rect 491 -30 503 30
rect 445 -42 503 -30
<< ndiffc >>
rect -491 -30 -457 30
rect -333 -30 -299 30
rect -175 -30 -141 30
rect -17 -30 17 30
rect 141 -30 175 30
rect 299 -30 333 30
rect 457 -30 491 30
<< psubdiff >>
rect -605 182 -509 216
rect 509 182 605 216
rect -605 120 -571 182
rect 571 120 605 182
rect -605 -182 -571 -120
rect 571 -182 605 -120
rect -605 -216 -509 -182
rect 509 -216 605 -182
<< psubdiffcont >>
rect -509 182 509 216
rect -605 -120 -571 120
rect 571 -120 605 120
rect -509 -216 509 -182
<< poly >>
rect -445 114 -345 130
rect -445 80 -429 114
rect -361 80 -345 114
rect -445 42 -345 80
rect -287 114 -187 130
rect -287 80 -271 114
rect -203 80 -187 114
rect -287 42 -187 80
rect -129 114 -29 130
rect -129 80 -113 114
rect -45 80 -29 114
rect -129 42 -29 80
rect 29 114 129 130
rect 29 80 45 114
rect 113 80 129 114
rect 29 42 129 80
rect 187 114 287 130
rect 187 80 203 114
rect 271 80 287 114
rect 187 42 287 80
rect 345 114 445 130
rect 345 80 361 114
rect 429 80 445 114
rect 345 42 445 80
rect -445 -80 -345 -42
rect -445 -114 -429 -80
rect -361 -114 -345 -80
rect -445 -130 -345 -114
rect -287 -80 -187 -42
rect -287 -114 -271 -80
rect -203 -114 -187 -80
rect -287 -130 -187 -114
rect -129 -80 -29 -42
rect -129 -114 -113 -80
rect -45 -114 -29 -80
rect -129 -130 -29 -114
rect 29 -80 129 -42
rect 29 -114 45 -80
rect 113 -114 129 -80
rect 29 -130 129 -114
rect 187 -80 287 -42
rect 187 -114 203 -80
rect 271 -114 287 -80
rect 187 -130 287 -114
rect 345 -80 445 -42
rect 345 -114 361 -80
rect 429 -114 445 -80
rect 345 -130 445 -114
<< polycont >>
rect -429 80 -361 114
rect -271 80 -203 114
rect -113 80 -45 114
rect 45 80 113 114
rect 203 80 271 114
rect 361 80 429 114
rect -429 -114 -361 -80
rect -271 -114 -203 -80
rect -113 -114 -45 -80
rect 45 -114 113 -80
rect 203 -114 271 -80
rect 361 -114 429 -80
<< locali >>
rect -605 182 -509 216
rect 509 182 605 216
rect -605 120 -571 182
rect 571 120 605 182
rect -445 80 -429 114
rect -361 80 -345 114
rect -287 80 -271 114
rect -203 80 -187 114
rect -129 80 -113 114
rect -45 80 -29 114
rect 29 80 45 114
rect 113 80 129 114
rect 187 80 203 114
rect 271 80 287 114
rect 345 80 361 114
rect 429 80 445 114
rect -491 30 -457 46
rect -491 -46 -457 -30
rect -333 30 -299 46
rect -333 -46 -299 -30
rect -175 30 -141 46
rect -175 -46 -141 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 141 30 175 46
rect 141 -46 175 -30
rect 299 30 333 46
rect 299 -46 333 -30
rect 457 30 491 46
rect 457 -46 491 -30
rect -445 -114 -429 -80
rect -361 -114 -345 -80
rect -287 -114 -271 -80
rect -203 -114 -187 -80
rect -129 -114 -113 -80
rect -45 -114 -29 -80
rect 29 -114 45 -80
rect 113 -114 129 -80
rect 187 -114 203 -80
rect 271 -114 287 -80
rect 345 -114 361 -80
rect 429 -114 445 -80
rect -605 -182 -571 -120
rect 571 -182 605 -120
rect -605 -216 -509 -182
rect 509 -216 605 -182
<< viali >>
rect -429 80 -361 114
rect -271 80 -203 114
rect -113 80 -45 114
rect 45 80 113 114
rect 203 80 271 114
rect 361 80 429 114
rect -491 -30 -457 30
rect -333 -30 -299 30
rect -175 -30 -141 30
rect -17 -30 17 30
rect 141 -30 175 30
rect 299 -30 333 30
rect 457 -30 491 30
rect -429 -114 -361 -80
rect -271 -114 -203 -80
rect -113 -114 -45 -80
rect 45 -114 113 -80
rect 203 -114 271 -80
rect 361 -114 429 -80
<< metal1 >>
rect -441 114 -349 120
rect -441 80 -429 114
rect -361 80 -349 114
rect -441 74 -349 80
rect -283 114 -191 120
rect -283 80 -271 114
rect -203 80 -191 114
rect -283 74 -191 80
rect -125 114 -33 120
rect -125 80 -113 114
rect -45 80 -33 114
rect -125 74 -33 80
rect 33 114 125 120
rect 33 80 45 114
rect 113 80 125 114
rect 33 74 125 80
rect 191 114 283 120
rect 191 80 203 114
rect 271 80 283 114
rect 191 74 283 80
rect 349 114 441 120
rect 349 80 361 114
rect 429 80 441 114
rect 349 74 441 80
rect -497 30 -451 42
rect -497 -30 -491 30
rect -457 -30 -451 30
rect -497 -42 -451 -30
rect -339 30 -293 42
rect -339 -30 -333 30
rect -299 -30 -293 30
rect -339 -42 -293 -30
rect -181 30 -135 42
rect -181 -30 -175 30
rect -141 -30 -135 30
rect -181 -42 -135 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 135 30 181 42
rect 135 -30 141 30
rect 175 -30 181 30
rect 135 -42 181 -30
rect 293 30 339 42
rect 293 -30 299 30
rect 333 -30 339 30
rect 293 -42 339 -30
rect 451 30 497 42
rect 451 -30 457 30
rect 491 -30 497 30
rect 451 -42 497 -30
rect -441 -80 -349 -74
rect -441 -114 -429 -80
rect -361 -114 -349 -80
rect -441 -120 -349 -114
rect -283 -80 -191 -74
rect -283 -114 -271 -80
rect -203 -114 -191 -80
rect -283 -120 -191 -114
rect -125 -80 -33 -74
rect -125 -114 -113 -80
rect -45 -114 -33 -80
rect -125 -120 -33 -114
rect 33 -80 125 -74
rect 33 -114 45 -80
rect 113 -114 125 -80
rect 33 -120 125 -114
rect 191 -80 283 -74
rect 191 -114 203 -80
rect 271 -114 283 -80
rect 191 -120 283 -114
rect 349 -80 441 -74
rect 349 -114 361 -80
rect 429 -114 441 -80
rect 349 -120 441 -114
<< properties >>
string FIXED_BBOX -588 -199 588 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.5 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
