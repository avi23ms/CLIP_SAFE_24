magic
tech sky130A
magscale 1 2
timestamp 1698317566
<< metal3 >>
rect 32 148 256 150
rect -86 -649 256 148
rect -90 -15462 261 -649
use capacitor_7  capacitor_7_0
timestamp 1698317566
transform 1 0 -9400 0 1 -938
box -32 0 9486 2050
use capacitor_7  capacitor_7_1
timestamp 1698317566
transform 1 0 -9400 0 1 -3022
box -32 0 9486 2050
use capacitor_7  capacitor_7_2
timestamp 1698317566
transform 1 0 -9408 0 1 -5106
box -32 0 9486 2050
use capacitor_7  capacitor_7_3
timestamp 1698317566
transform 1 0 -9414 0 1 -7190
box -32 0 9486 2050
use capacitor_7  capacitor_7_4
timestamp 1698317566
transform 1 0 -9400 0 1 -9272
box -32 0 9486 2050
use capacitor_7  capacitor_7_5
timestamp 1698317566
transform 1 0 -9400 0 1 -11356
box -32 0 9486 2050
use capacitor_7  capacitor_7_6
timestamp 1698317566
transform 1 0 -9400 0 1 -13440
box -32 0 9486 2050
use capacitor_7  capacitor_7_7
timestamp 1698317566
transform 1 0 -9400 0 1 -15524
box -32 0 9486 2050
<< end >>
