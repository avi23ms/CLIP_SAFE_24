magic
tech sky130A
magscale 1 2
timestamp 1698659501
<< nmos >>
rect -2847 -42 -2817 42
rect -2751 -42 -2721 42
rect -2655 -42 -2625 42
rect -2559 -42 -2529 42
rect -2463 -42 -2433 42
rect -2367 -42 -2337 42
rect -2271 -42 -2241 42
rect -2175 -42 -2145 42
rect -2079 -42 -2049 42
rect -1983 -42 -1953 42
rect -1887 -42 -1857 42
rect -1791 -42 -1761 42
rect -1695 -42 -1665 42
rect -1599 -42 -1569 42
rect -1503 -42 -1473 42
rect -1407 -42 -1377 42
rect -1311 -42 -1281 42
rect -1215 -42 -1185 42
rect -1119 -42 -1089 42
rect -1023 -42 -993 42
rect -927 -42 -897 42
rect -831 -42 -801 42
rect -735 -42 -705 42
rect -639 -42 -609 42
rect -543 -42 -513 42
rect -447 -42 -417 42
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
rect 417 -42 447 42
rect 513 -42 543 42
rect 609 -42 639 42
rect 705 -42 735 42
rect 801 -42 831 42
rect 897 -42 927 42
rect 993 -42 1023 42
rect 1089 -42 1119 42
rect 1185 -42 1215 42
rect 1281 -42 1311 42
rect 1377 -42 1407 42
rect 1473 -42 1503 42
rect 1569 -42 1599 42
rect 1665 -42 1695 42
rect 1761 -42 1791 42
rect 1857 -42 1887 42
rect 1953 -42 1983 42
rect 2049 -42 2079 42
rect 2145 -42 2175 42
rect 2241 -42 2271 42
rect 2337 -42 2367 42
rect 2433 -42 2463 42
rect 2529 -42 2559 42
rect 2625 -42 2655 42
rect 2721 -42 2751 42
rect 2817 -42 2847 42
<< ndiff >>
rect -2909 30 -2847 42
rect -2909 -30 -2897 30
rect -2863 -30 -2847 30
rect -2909 -42 -2847 -30
rect -2817 30 -2751 42
rect -2817 -30 -2801 30
rect -2767 -30 -2751 30
rect -2817 -42 -2751 -30
rect -2721 30 -2655 42
rect -2721 -30 -2705 30
rect -2671 -30 -2655 30
rect -2721 -42 -2655 -30
rect -2625 30 -2559 42
rect -2625 -30 -2609 30
rect -2575 -30 -2559 30
rect -2625 -42 -2559 -30
rect -2529 30 -2463 42
rect -2529 -30 -2513 30
rect -2479 -30 -2463 30
rect -2529 -42 -2463 -30
rect -2433 30 -2367 42
rect -2433 -30 -2417 30
rect -2383 -30 -2367 30
rect -2433 -42 -2367 -30
rect -2337 30 -2271 42
rect -2337 -30 -2321 30
rect -2287 -30 -2271 30
rect -2337 -42 -2271 -30
rect -2241 30 -2175 42
rect -2241 -30 -2225 30
rect -2191 -30 -2175 30
rect -2241 -42 -2175 -30
rect -2145 30 -2079 42
rect -2145 -30 -2129 30
rect -2095 -30 -2079 30
rect -2145 -42 -2079 -30
rect -2049 30 -1983 42
rect -2049 -30 -2033 30
rect -1999 -30 -1983 30
rect -2049 -42 -1983 -30
rect -1953 30 -1887 42
rect -1953 -30 -1937 30
rect -1903 -30 -1887 30
rect -1953 -42 -1887 -30
rect -1857 30 -1791 42
rect -1857 -30 -1841 30
rect -1807 -30 -1791 30
rect -1857 -42 -1791 -30
rect -1761 30 -1695 42
rect -1761 -30 -1745 30
rect -1711 -30 -1695 30
rect -1761 -42 -1695 -30
rect -1665 30 -1599 42
rect -1665 -30 -1649 30
rect -1615 -30 -1599 30
rect -1665 -42 -1599 -30
rect -1569 30 -1503 42
rect -1569 -30 -1553 30
rect -1519 -30 -1503 30
rect -1569 -42 -1503 -30
rect -1473 30 -1407 42
rect -1473 -30 -1457 30
rect -1423 -30 -1407 30
rect -1473 -42 -1407 -30
rect -1377 30 -1311 42
rect -1377 -30 -1361 30
rect -1327 -30 -1311 30
rect -1377 -42 -1311 -30
rect -1281 30 -1215 42
rect -1281 -30 -1265 30
rect -1231 -30 -1215 30
rect -1281 -42 -1215 -30
rect -1185 30 -1119 42
rect -1185 -30 -1169 30
rect -1135 -30 -1119 30
rect -1185 -42 -1119 -30
rect -1089 30 -1023 42
rect -1089 -30 -1073 30
rect -1039 -30 -1023 30
rect -1089 -42 -1023 -30
rect -993 30 -927 42
rect -993 -30 -977 30
rect -943 -30 -927 30
rect -993 -42 -927 -30
rect -897 30 -831 42
rect -897 -30 -881 30
rect -847 -30 -831 30
rect -897 -42 -831 -30
rect -801 30 -735 42
rect -801 -30 -785 30
rect -751 -30 -735 30
rect -801 -42 -735 -30
rect -705 30 -639 42
rect -705 -30 -689 30
rect -655 -30 -639 30
rect -705 -42 -639 -30
rect -609 30 -543 42
rect -609 -30 -593 30
rect -559 -30 -543 30
rect -609 -42 -543 -30
rect -513 30 -447 42
rect -513 -30 -497 30
rect -463 -30 -447 30
rect -513 -42 -447 -30
rect -417 30 -351 42
rect -417 -30 -401 30
rect -367 -30 -351 30
rect -417 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 417 42
rect 351 -30 367 30
rect 401 -30 417 30
rect 351 -42 417 -30
rect 447 30 513 42
rect 447 -30 463 30
rect 497 -30 513 30
rect 447 -42 513 -30
rect 543 30 609 42
rect 543 -30 559 30
rect 593 -30 609 30
rect 543 -42 609 -30
rect 639 30 705 42
rect 639 -30 655 30
rect 689 -30 705 30
rect 639 -42 705 -30
rect 735 30 801 42
rect 735 -30 751 30
rect 785 -30 801 30
rect 735 -42 801 -30
rect 831 30 897 42
rect 831 -30 847 30
rect 881 -30 897 30
rect 831 -42 897 -30
rect 927 30 993 42
rect 927 -30 943 30
rect 977 -30 993 30
rect 927 -42 993 -30
rect 1023 30 1089 42
rect 1023 -30 1039 30
rect 1073 -30 1089 30
rect 1023 -42 1089 -30
rect 1119 30 1185 42
rect 1119 -30 1135 30
rect 1169 -30 1185 30
rect 1119 -42 1185 -30
rect 1215 30 1281 42
rect 1215 -30 1231 30
rect 1265 -30 1281 30
rect 1215 -42 1281 -30
rect 1311 30 1377 42
rect 1311 -30 1327 30
rect 1361 -30 1377 30
rect 1311 -42 1377 -30
rect 1407 30 1473 42
rect 1407 -30 1423 30
rect 1457 -30 1473 30
rect 1407 -42 1473 -30
rect 1503 30 1569 42
rect 1503 -30 1519 30
rect 1553 -30 1569 30
rect 1503 -42 1569 -30
rect 1599 30 1665 42
rect 1599 -30 1615 30
rect 1649 -30 1665 30
rect 1599 -42 1665 -30
rect 1695 30 1761 42
rect 1695 -30 1711 30
rect 1745 -30 1761 30
rect 1695 -42 1761 -30
rect 1791 30 1857 42
rect 1791 -30 1807 30
rect 1841 -30 1857 30
rect 1791 -42 1857 -30
rect 1887 30 1953 42
rect 1887 -30 1903 30
rect 1937 -30 1953 30
rect 1887 -42 1953 -30
rect 1983 30 2049 42
rect 1983 -30 1999 30
rect 2033 -30 2049 30
rect 1983 -42 2049 -30
rect 2079 30 2145 42
rect 2079 -30 2095 30
rect 2129 -30 2145 30
rect 2079 -42 2145 -30
rect 2175 30 2241 42
rect 2175 -30 2191 30
rect 2225 -30 2241 30
rect 2175 -42 2241 -30
rect 2271 30 2337 42
rect 2271 -30 2287 30
rect 2321 -30 2337 30
rect 2271 -42 2337 -30
rect 2367 30 2433 42
rect 2367 -30 2383 30
rect 2417 -30 2433 30
rect 2367 -42 2433 -30
rect 2463 30 2529 42
rect 2463 -30 2479 30
rect 2513 -30 2529 30
rect 2463 -42 2529 -30
rect 2559 30 2625 42
rect 2559 -30 2575 30
rect 2609 -30 2625 30
rect 2559 -42 2625 -30
rect 2655 30 2721 42
rect 2655 -30 2671 30
rect 2705 -30 2721 30
rect 2655 -42 2721 -30
rect 2751 30 2817 42
rect 2751 -30 2767 30
rect 2801 -30 2817 30
rect 2751 -42 2817 -30
rect 2847 30 2909 42
rect 2847 -30 2863 30
rect 2897 -30 2909 30
rect 2847 -42 2909 -30
<< ndiffc >>
rect -2897 -30 -2863 30
rect -2801 -30 -2767 30
rect -2705 -30 -2671 30
rect -2609 -30 -2575 30
rect -2513 -30 -2479 30
rect -2417 -30 -2383 30
rect -2321 -30 -2287 30
rect -2225 -30 -2191 30
rect -2129 -30 -2095 30
rect -2033 -30 -1999 30
rect -1937 -30 -1903 30
rect -1841 -30 -1807 30
rect -1745 -30 -1711 30
rect -1649 -30 -1615 30
rect -1553 -30 -1519 30
rect -1457 -30 -1423 30
rect -1361 -30 -1327 30
rect -1265 -30 -1231 30
rect -1169 -30 -1135 30
rect -1073 -30 -1039 30
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
rect 1039 -30 1073 30
rect 1135 -30 1169 30
rect 1231 -30 1265 30
rect 1327 -30 1361 30
rect 1423 -30 1457 30
rect 1519 -30 1553 30
rect 1615 -30 1649 30
rect 1711 -30 1745 30
rect 1807 -30 1841 30
rect 1903 -30 1937 30
rect 1999 -30 2033 30
rect 2095 -30 2129 30
rect 2191 -30 2225 30
rect 2287 -30 2321 30
rect 2383 -30 2417 30
rect 2479 -30 2513 30
rect 2575 -30 2609 30
rect 2671 -30 2705 30
rect 2767 -30 2801 30
rect 2863 -30 2897 30
<< poly >>
rect -2769 114 -2703 130
rect -2769 80 -2753 114
rect -2719 80 -2703 114
rect -2847 42 -2817 68
rect -2769 64 -2703 80
rect -2577 114 -2511 130
rect -2577 80 -2561 114
rect -2527 80 -2511 114
rect -2751 42 -2721 64
rect -2655 42 -2625 68
rect -2577 64 -2511 80
rect -2385 114 -2319 130
rect -2385 80 -2369 114
rect -2335 80 -2319 114
rect -2559 42 -2529 64
rect -2463 42 -2433 68
rect -2385 64 -2319 80
rect -2193 114 -2127 130
rect -2193 80 -2177 114
rect -2143 80 -2127 114
rect -2367 42 -2337 64
rect -2271 42 -2241 68
rect -2193 64 -2127 80
rect -2001 114 -1935 130
rect -2001 80 -1985 114
rect -1951 80 -1935 114
rect -2175 42 -2145 64
rect -2079 42 -2049 68
rect -2001 64 -1935 80
rect -1809 114 -1743 130
rect -1809 80 -1793 114
rect -1759 80 -1743 114
rect -1983 42 -1953 64
rect -1887 42 -1857 68
rect -1809 64 -1743 80
rect -1617 114 -1551 130
rect -1617 80 -1601 114
rect -1567 80 -1551 114
rect -1791 42 -1761 64
rect -1695 42 -1665 68
rect -1617 64 -1551 80
rect -1425 114 -1359 130
rect -1425 80 -1409 114
rect -1375 80 -1359 114
rect -1599 42 -1569 64
rect -1503 42 -1473 68
rect -1425 64 -1359 80
rect -1233 114 -1167 130
rect -1233 80 -1217 114
rect -1183 80 -1167 114
rect -1407 42 -1377 64
rect -1311 42 -1281 68
rect -1233 64 -1167 80
rect -1041 114 -975 130
rect -1041 80 -1025 114
rect -991 80 -975 114
rect -1215 42 -1185 64
rect -1119 42 -1089 68
rect -1041 64 -975 80
rect -849 114 -783 130
rect -849 80 -833 114
rect -799 80 -783 114
rect -1023 42 -993 64
rect -927 42 -897 68
rect -849 64 -783 80
rect -657 114 -591 130
rect -657 80 -641 114
rect -607 80 -591 114
rect -831 42 -801 64
rect -735 42 -705 68
rect -657 64 -591 80
rect -465 114 -399 130
rect -465 80 -449 114
rect -415 80 -399 114
rect -639 42 -609 64
rect -543 42 -513 68
rect -465 64 -399 80
rect -273 114 -207 130
rect -273 80 -257 114
rect -223 80 -207 114
rect -447 42 -417 64
rect -351 42 -321 68
rect -273 64 -207 80
rect -81 114 -15 130
rect -81 80 -65 114
rect -31 80 -15 114
rect -255 42 -225 64
rect -159 42 -129 68
rect -81 64 -15 80
rect 111 114 177 130
rect 111 80 127 114
rect 161 80 177 114
rect -63 42 -33 64
rect 33 42 63 68
rect 111 64 177 80
rect 303 114 369 130
rect 303 80 319 114
rect 353 80 369 114
rect 129 42 159 64
rect 225 42 255 68
rect 303 64 369 80
rect 495 114 561 130
rect 495 80 511 114
rect 545 80 561 114
rect 321 42 351 64
rect 417 42 447 68
rect 495 64 561 80
rect 687 114 753 130
rect 687 80 703 114
rect 737 80 753 114
rect 513 42 543 64
rect 609 42 639 68
rect 687 64 753 80
rect 879 114 945 130
rect 879 80 895 114
rect 929 80 945 114
rect 705 42 735 64
rect 801 42 831 68
rect 879 64 945 80
rect 1071 114 1137 130
rect 1071 80 1087 114
rect 1121 80 1137 114
rect 897 42 927 64
rect 993 42 1023 68
rect 1071 64 1137 80
rect 1263 114 1329 130
rect 1263 80 1279 114
rect 1313 80 1329 114
rect 1089 42 1119 64
rect 1185 42 1215 68
rect 1263 64 1329 80
rect 1455 114 1521 130
rect 1455 80 1471 114
rect 1505 80 1521 114
rect 1281 42 1311 64
rect 1377 42 1407 68
rect 1455 64 1521 80
rect 1647 114 1713 130
rect 1647 80 1663 114
rect 1697 80 1713 114
rect 1473 42 1503 64
rect 1569 42 1599 68
rect 1647 64 1713 80
rect 1839 114 1905 130
rect 1839 80 1855 114
rect 1889 80 1905 114
rect 1665 42 1695 64
rect 1761 42 1791 68
rect 1839 64 1905 80
rect 2031 114 2097 130
rect 2031 80 2047 114
rect 2081 80 2097 114
rect 1857 42 1887 64
rect 1953 42 1983 68
rect 2031 64 2097 80
rect 2223 114 2289 130
rect 2223 80 2239 114
rect 2273 80 2289 114
rect 2049 42 2079 64
rect 2145 42 2175 68
rect 2223 64 2289 80
rect 2415 114 2481 130
rect 2415 80 2431 114
rect 2465 80 2481 114
rect 2241 42 2271 64
rect 2337 42 2367 68
rect 2415 64 2481 80
rect 2607 114 2673 130
rect 2607 80 2623 114
rect 2657 80 2673 114
rect 2433 42 2463 64
rect 2529 42 2559 68
rect 2607 64 2673 80
rect 2799 114 2865 130
rect 2799 80 2815 114
rect 2849 80 2865 114
rect 2625 42 2655 64
rect 2721 42 2751 68
rect 2799 64 2865 80
rect 2817 42 2847 64
rect -2847 -64 -2817 -42
rect -2865 -80 -2799 -64
rect -2751 -68 -2721 -42
rect -2655 -64 -2625 -42
rect -2865 -114 -2849 -80
rect -2815 -114 -2799 -80
rect -2865 -130 -2799 -114
rect -2673 -80 -2607 -64
rect -2559 -68 -2529 -42
rect -2463 -64 -2433 -42
rect -2673 -114 -2657 -80
rect -2623 -114 -2607 -80
rect -2673 -130 -2607 -114
rect -2481 -80 -2415 -64
rect -2367 -68 -2337 -42
rect -2271 -64 -2241 -42
rect -2481 -114 -2465 -80
rect -2431 -114 -2415 -80
rect -2481 -130 -2415 -114
rect -2289 -80 -2223 -64
rect -2175 -68 -2145 -42
rect -2079 -64 -2049 -42
rect -2289 -114 -2273 -80
rect -2239 -114 -2223 -80
rect -2289 -130 -2223 -114
rect -2097 -80 -2031 -64
rect -1983 -68 -1953 -42
rect -1887 -64 -1857 -42
rect -2097 -114 -2081 -80
rect -2047 -114 -2031 -80
rect -2097 -130 -2031 -114
rect -1905 -80 -1839 -64
rect -1791 -68 -1761 -42
rect -1695 -64 -1665 -42
rect -1905 -114 -1889 -80
rect -1855 -114 -1839 -80
rect -1905 -130 -1839 -114
rect -1713 -80 -1647 -64
rect -1599 -68 -1569 -42
rect -1503 -64 -1473 -42
rect -1713 -114 -1697 -80
rect -1663 -114 -1647 -80
rect -1713 -130 -1647 -114
rect -1521 -80 -1455 -64
rect -1407 -68 -1377 -42
rect -1311 -64 -1281 -42
rect -1521 -114 -1505 -80
rect -1471 -114 -1455 -80
rect -1521 -130 -1455 -114
rect -1329 -80 -1263 -64
rect -1215 -68 -1185 -42
rect -1119 -64 -1089 -42
rect -1329 -114 -1313 -80
rect -1279 -114 -1263 -80
rect -1329 -130 -1263 -114
rect -1137 -80 -1071 -64
rect -1023 -68 -993 -42
rect -927 -64 -897 -42
rect -1137 -114 -1121 -80
rect -1087 -114 -1071 -80
rect -1137 -130 -1071 -114
rect -945 -80 -879 -64
rect -831 -68 -801 -42
rect -735 -64 -705 -42
rect -945 -114 -929 -80
rect -895 -114 -879 -80
rect -945 -130 -879 -114
rect -753 -80 -687 -64
rect -639 -68 -609 -42
rect -543 -64 -513 -42
rect -753 -114 -737 -80
rect -703 -114 -687 -80
rect -753 -130 -687 -114
rect -561 -80 -495 -64
rect -447 -68 -417 -42
rect -351 -64 -321 -42
rect -561 -114 -545 -80
rect -511 -114 -495 -80
rect -561 -130 -495 -114
rect -369 -80 -303 -64
rect -255 -68 -225 -42
rect -159 -64 -129 -42
rect -369 -114 -353 -80
rect -319 -114 -303 -80
rect -369 -130 -303 -114
rect -177 -80 -111 -64
rect -63 -68 -33 -42
rect 33 -64 63 -42
rect -177 -114 -161 -80
rect -127 -114 -111 -80
rect -177 -130 -111 -114
rect 15 -80 81 -64
rect 129 -68 159 -42
rect 225 -64 255 -42
rect 15 -114 31 -80
rect 65 -114 81 -80
rect 15 -130 81 -114
rect 207 -80 273 -64
rect 321 -68 351 -42
rect 417 -64 447 -42
rect 207 -114 223 -80
rect 257 -114 273 -80
rect 207 -130 273 -114
rect 399 -80 465 -64
rect 513 -68 543 -42
rect 609 -64 639 -42
rect 399 -114 415 -80
rect 449 -114 465 -80
rect 399 -130 465 -114
rect 591 -80 657 -64
rect 705 -68 735 -42
rect 801 -64 831 -42
rect 591 -114 607 -80
rect 641 -114 657 -80
rect 591 -130 657 -114
rect 783 -80 849 -64
rect 897 -68 927 -42
rect 993 -64 1023 -42
rect 783 -114 799 -80
rect 833 -114 849 -80
rect 783 -130 849 -114
rect 975 -80 1041 -64
rect 1089 -68 1119 -42
rect 1185 -64 1215 -42
rect 975 -114 991 -80
rect 1025 -114 1041 -80
rect 975 -130 1041 -114
rect 1167 -80 1233 -64
rect 1281 -68 1311 -42
rect 1377 -64 1407 -42
rect 1167 -114 1183 -80
rect 1217 -114 1233 -80
rect 1167 -130 1233 -114
rect 1359 -80 1425 -64
rect 1473 -68 1503 -42
rect 1569 -64 1599 -42
rect 1359 -114 1375 -80
rect 1409 -114 1425 -80
rect 1359 -130 1425 -114
rect 1551 -80 1617 -64
rect 1665 -68 1695 -42
rect 1761 -64 1791 -42
rect 1551 -114 1567 -80
rect 1601 -114 1617 -80
rect 1551 -130 1617 -114
rect 1743 -80 1809 -64
rect 1857 -68 1887 -42
rect 1953 -64 1983 -42
rect 1743 -114 1759 -80
rect 1793 -114 1809 -80
rect 1743 -130 1809 -114
rect 1935 -80 2001 -64
rect 2049 -68 2079 -42
rect 2145 -64 2175 -42
rect 1935 -114 1951 -80
rect 1985 -114 2001 -80
rect 1935 -130 2001 -114
rect 2127 -80 2193 -64
rect 2241 -68 2271 -42
rect 2337 -64 2367 -42
rect 2127 -114 2143 -80
rect 2177 -114 2193 -80
rect 2127 -130 2193 -114
rect 2319 -80 2385 -64
rect 2433 -68 2463 -42
rect 2529 -64 2559 -42
rect 2319 -114 2335 -80
rect 2369 -114 2385 -80
rect 2319 -130 2385 -114
rect 2511 -80 2577 -64
rect 2625 -68 2655 -42
rect 2721 -64 2751 -42
rect 2511 -114 2527 -80
rect 2561 -114 2577 -80
rect 2511 -130 2577 -114
rect 2703 -80 2769 -64
rect 2817 -68 2847 -42
rect 2703 -114 2719 -80
rect 2753 -114 2769 -80
rect 2703 -130 2769 -114
<< polycont >>
rect -2753 80 -2719 114
rect -2561 80 -2527 114
rect -2369 80 -2335 114
rect -2177 80 -2143 114
rect -1985 80 -1951 114
rect -1793 80 -1759 114
rect -1601 80 -1567 114
rect -1409 80 -1375 114
rect -1217 80 -1183 114
rect -1025 80 -991 114
rect -833 80 -799 114
rect -641 80 -607 114
rect -449 80 -415 114
rect -257 80 -223 114
rect -65 80 -31 114
rect 127 80 161 114
rect 319 80 353 114
rect 511 80 545 114
rect 703 80 737 114
rect 895 80 929 114
rect 1087 80 1121 114
rect 1279 80 1313 114
rect 1471 80 1505 114
rect 1663 80 1697 114
rect 1855 80 1889 114
rect 2047 80 2081 114
rect 2239 80 2273 114
rect 2431 80 2465 114
rect 2623 80 2657 114
rect 2815 80 2849 114
rect -2849 -114 -2815 -80
rect -2657 -114 -2623 -80
rect -2465 -114 -2431 -80
rect -2273 -114 -2239 -80
rect -2081 -114 -2047 -80
rect -1889 -114 -1855 -80
rect -1697 -114 -1663 -80
rect -1505 -114 -1471 -80
rect -1313 -114 -1279 -80
rect -1121 -114 -1087 -80
rect -929 -114 -895 -80
rect -737 -114 -703 -80
rect -545 -114 -511 -80
rect -353 -114 -319 -80
rect -161 -114 -127 -80
rect 31 -114 65 -80
rect 223 -114 257 -80
rect 415 -114 449 -80
rect 607 -114 641 -80
rect 799 -114 833 -80
rect 991 -114 1025 -80
rect 1183 -114 1217 -80
rect 1375 -114 1409 -80
rect 1567 -114 1601 -80
rect 1759 -114 1793 -80
rect 1951 -114 1985 -80
rect 2143 -114 2177 -80
rect 2335 -114 2369 -80
rect 2527 -114 2561 -80
rect 2719 -114 2753 -80
<< locali >>
rect -2769 80 -2753 114
rect -2719 80 -2703 114
rect -2577 80 -2561 114
rect -2527 80 -2511 114
rect -2385 80 -2369 114
rect -2335 80 -2319 114
rect -2193 80 -2177 114
rect -2143 80 -2127 114
rect -2001 80 -1985 114
rect -1951 80 -1935 114
rect -1809 80 -1793 114
rect -1759 80 -1743 114
rect -1617 80 -1601 114
rect -1567 80 -1551 114
rect -1425 80 -1409 114
rect -1375 80 -1359 114
rect -1233 80 -1217 114
rect -1183 80 -1167 114
rect -1041 80 -1025 114
rect -991 80 -975 114
rect -849 80 -833 114
rect -799 80 -783 114
rect -657 80 -641 114
rect -607 80 -591 114
rect -465 80 -449 114
rect -415 80 -399 114
rect -273 80 -257 114
rect -223 80 -207 114
rect -81 80 -65 114
rect -31 80 -15 114
rect 111 80 127 114
rect 161 80 177 114
rect 303 80 319 114
rect 353 80 369 114
rect 495 80 511 114
rect 545 80 561 114
rect 687 80 703 114
rect 737 80 753 114
rect 879 80 895 114
rect 929 80 945 114
rect 1071 80 1087 114
rect 1121 80 1137 114
rect 1263 80 1279 114
rect 1313 80 1329 114
rect 1455 80 1471 114
rect 1505 80 1521 114
rect 1647 80 1663 114
rect 1697 80 1713 114
rect 1839 80 1855 114
rect 1889 80 1905 114
rect 2031 80 2047 114
rect 2081 80 2097 114
rect 2223 80 2239 114
rect 2273 80 2289 114
rect 2415 80 2431 114
rect 2465 80 2481 114
rect 2607 80 2623 114
rect 2657 80 2673 114
rect 2799 80 2815 114
rect 2849 80 2865 114
rect -2897 30 -2863 46
rect -2897 -46 -2863 -30
rect -2801 30 -2767 46
rect -2801 -46 -2767 -30
rect -2705 30 -2671 46
rect -2705 -46 -2671 -30
rect -2609 30 -2575 46
rect -2609 -46 -2575 -30
rect -2513 30 -2479 46
rect -2513 -46 -2479 -30
rect -2417 30 -2383 46
rect -2417 -46 -2383 -30
rect -2321 30 -2287 46
rect -2321 -46 -2287 -30
rect -2225 30 -2191 46
rect -2225 -46 -2191 -30
rect -2129 30 -2095 46
rect -2129 -46 -2095 -30
rect -2033 30 -1999 46
rect -2033 -46 -1999 -30
rect -1937 30 -1903 46
rect -1937 -46 -1903 -30
rect -1841 30 -1807 46
rect -1841 -46 -1807 -30
rect -1745 30 -1711 46
rect -1745 -46 -1711 -30
rect -1649 30 -1615 46
rect -1649 -46 -1615 -30
rect -1553 30 -1519 46
rect -1553 -46 -1519 -30
rect -1457 30 -1423 46
rect -1457 -46 -1423 -30
rect -1361 30 -1327 46
rect -1361 -46 -1327 -30
rect -1265 30 -1231 46
rect -1265 -46 -1231 -30
rect -1169 30 -1135 46
rect -1169 -46 -1135 -30
rect -1073 30 -1039 46
rect -1073 -46 -1039 -30
rect -977 30 -943 46
rect -977 -46 -943 -30
rect -881 30 -847 46
rect -881 -46 -847 -30
rect -785 30 -751 46
rect -785 -46 -751 -30
rect -689 30 -655 46
rect -689 -46 -655 -30
rect -593 30 -559 46
rect -593 -46 -559 -30
rect -497 30 -463 46
rect -497 -46 -463 -30
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect 463 30 497 46
rect 463 -46 497 -30
rect 559 30 593 46
rect 559 -46 593 -30
rect 655 30 689 46
rect 655 -46 689 -30
rect 751 30 785 46
rect 751 -46 785 -30
rect 847 30 881 46
rect 847 -46 881 -30
rect 943 30 977 46
rect 943 -46 977 -30
rect 1039 30 1073 46
rect 1039 -46 1073 -30
rect 1135 30 1169 46
rect 1135 -46 1169 -30
rect 1231 30 1265 46
rect 1231 -46 1265 -30
rect 1327 30 1361 46
rect 1327 -46 1361 -30
rect 1423 30 1457 46
rect 1423 -46 1457 -30
rect 1519 30 1553 46
rect 1519 -46 1553 -30
rect 1615 30 1649 46
rect 1615 -46 1649 -30
rect 1711 30 1745 46
rect 1711 -46 1745 -30
rect 1807 30 1841 46
rect 1807 -46 1841 -30
rect 1903 30 1937 46
rect 1903 -46 1937 -30
rect 1999 30 2033 46
rect 1999 -46 2033 -30
rect 2095 30 2129 46
rect 2095 -46 2129 -30
rect 2191 30 2225 46
rect 2191 -46 2225 -30
rect 2287 30 2321 46
rect 2287 -46 2321 -30
rect 2383 30 2417 46
rect 2383 -46 2417 -30
rect 2479 30 2513 46
rect 2479 -46 2513 -30
rect 2575 30 2609 46
rect 2575 -46 2609 -30
rect 2671 30 2705 46
rect 2671 -46 2705 -30
rect 2767 30 2801 46
rect 2767 -46 2801 -30
rect 2863 30 2897 46
rect 2863 -46 2897 -30
rect -2865 -114 -2849 -80
rect -2815 -114 -2799 -80
rect -2673 -114 -2657 -80
rect -2623 -114 -2607 -80
rect -2481 -114 -2465 -80
rect -2431 -114 -2415 -80
rect -2289 -114 -2273 -80
rect -2239 -114 -2223 -80
rect -2097 -114 -2081 -80
rect -2047 -114 -2031 -80
rect -1905 -114 -1889 -80
rect -1855 -114 -1839 -80
rect -1713 -114 -1697 -80
rect -1663 -114 -1647 -80
rect -1521 -114 -1505 -80
rect -1471 -114 -1455 -80
rect -1329 -114 -1313 -80
rect -1279 -114 -1263 -80
rect -1137 -114 -1121 -80
rect -1087 -114 -1071 -80
rect -945 -114 -929 -80
rect -895 -114 -879 -80
rect -753 -114 -737 -80
rect -703 -114 -687 -80
rect -561 -114 -545 -80
rect -511 -114 -495 -80
rect -369 -114 -353 -80
rect -319 -114 -303 -80
rect -177 -114 -161 -80
rect -127 -114 -111 -80
rect 15 -114 31 -80
rect 65 -114 81 -80
rect 207 -114 223 -80
rect 257 -114 273 -80
rect 399 -114 415 -80
rect 449 -114 465 -80
rect 591 -114 607 -80
rect 641 -114 657 -80
rect 783 -114 799 -80
rect 833 -114 849 -80
rect 975 -114 991 -80
rect 1025 -114 1041 -80
rect 1167 -114 1183 -80
rect 1217 -114 1233 -80
rect 1359 -114 1375 -80
rect 1409 -114 1425 -80
rect 1551 -114 1567 -80
rect 1601 -114 1617 -80
rect 1743 -114 1759 -80
rect 1793 -114 1809 -80
rect 1935 -114 1951 -80
rect 1985 -114 2001 -80
rect 2127 -114 2143 -80
rect 2177 -114 2193 -80
rect 2319 -114 2335 -80
rect 2369 -114 2385 -80
rect 2511 -114 2527 -80
rect 2561 -114 2577 -80
rect 2703 -114 2719 -80
rect 2753 -114 2769 -80
<< viali >>
rect -2897 -30 -2863 30
rect -2801 -30 -2767 30
rect -2705 -30 -2671 30
rect -2609 -30 -2575 30
rect -2513 -30 -2479 30
rect -2417 -30 -2383 30
rect -2321 -30 -2287 30
rect -2225 -30 -2191 30
rect -2129 -30 -2095 30
rect -2033 -30 -1999 30
rect -1937 -30 -1903 30
rect -1841 -30 -1807 30
rect -1745 -30 -1711 30
rect -1649 -30 -1615 30
rect -1553 -30 -1519 30
rect -1457 -30 -1423 30
rect -1361 -30 -1327 30
rect -1265 -30 -1231 30
rect -1169 -30 -1135 30
rect -1073 -30 -1039 30
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
rect 1039 -30 1073 30
rect 1135 -30 1169 30
rect 1231 -30 1265 30
rect 1327 -30 1361 30
rect 1423 -30 1457 30
rect 1519 -30 1553 30
rect 1615 -30 1649 30
rect 1711 -30 1745 30
rect 1807 -30 1841 30
rect 1903 -30 1937 30
rect 1999 -30 2033 30
rect 2095 -30 2129 30
rect 2191 -30 2225 30
rect 2287 -30 2321 30
rect 2383 -30 2417 30
rect 2479 -30 2513 30
rect 2575 -30 2609 30
rect 2671 -30 2705 30
rect 2767 -30 2801 30
rect 2863 -30 2897 30
<< metal1 >>
rect -2903 30 -2857 42
rect -2903 -30 -2897 30
rect -2863 -30 -2857 30
rect -2903 -42 -2857 -30
rect -2807 30 -2761 42
rect -2807 -30 -2801 30
rect -2767 -30 -2761 30
rect -2807 -42 -2761 -30
rect -2711 30 -2665 42
rect -2711 -30 -2705 30
rect -2671 -30 -2665 30
rect -2711 -42 -2665 -30
rect -2615 30 -2569 42
rect -2615 -30 -2609 30
rect -2575 -30 -2569 30
rect -2615 -42 -2569 -30
rect -2519 30 -2473 42
rect -2519 -30 -2513 30
rect -2479 -30 -2473 30
rect -2519 -42 -2473 -30
rect -2423 30 -2377 42
rect -2423 -30 -2417 30
rect -2383 -30 -2377 30
rect -2423 -42 -2377 -30
rect -2327 30 -2281 42
rect -2327 -30 -2321 30
rect -2287 -30 -2281 30
rect -2327 -42 -2281 -30
rect -2231 30 -2185 42
rect -2231 -30 -2225 30
rect -2191 -30 -2185 30
rect -2231 -42 -2185 -30
rect -2135 30 -2089 42
rect -2135 -30 -2129 30
rect -2095 -30 -2089 30
rect -2135 -42 -2089 -30
rect -2039 30 -1993 42
rect -2039 -30 -2033 30
rect -1999 -30 -1993 30
rect -2039 -42 -1993 -30
rect -1943 30 -1897 42
rect -1943 -30 -1937 30
rect -1903 -30 -1897 30
rect -1943 -42 -1897 -30
rect -1847 30 -1801 42
rect -1847 -30 -1841 30
rect -1807 -30 -1801 30
rect -1847 -42 -1801 -30
rect -1751 30 -1705 42
rect -1751 -30 -1745 30
rect -1711 -30 -1705 30
rect -1751 -42 -1705 -30
rect -1655 30 -1609 42
rect -1655 -30 -1649 30
rect -1615 -30 -1609 30
rect -1655 -42 -1609 -30
rect -1559 30 -1513 42
rect -1559 -30 -1553 30
rect -1519 -30 -1513 30
rect -1559 -42 -1513 -30
rect -1463 30 -1417 42
rect -1463 -30 -1457 30
rect -1423 -30 -1417 30
rect -1463 -42 -1417 -30
rect -1367 30 -1321 42
rect -1367 -30 -1361 30
rect -1327 -30 -1321 30
rect -1367 -42 -1321 -30
rect -1271 30 -1225 42
rect -1271 -30 -1265 30
rect -1231 -30 -1225 30
rect -1271 -42 -1225 -30
rect -1175 30 -1129 42
rect -1175 -30 -1169 30
rect -1135 -30 -1129 30
rect -1175 -42 -1129 -30
rect -1079 30 -1033 42
rect -1079 -30 -1073 30
rect -1039 -30 -1033 30
rect -1079 -42 -1033 -30
rect -983 30 -937 42
rect -983 -30 -977 30
rect -943 -30 -937 30
rect -983 -42 -937 -30
rect -887 30 -841 42
rect -887 -30 -881 30
rect -847 -30 -841 30
rect -887 -42 -841 -30
rect -791 30 -745 42
rect -791 -30 -785 30
rect -751 -30 -745 30
rect -791 -42 -745 -30
rect -695 30 -649 42
rect -695 -30 -689 30
rect -655 -30 -649 30
rect -695 -42 -649 -30
rect -599 30 -553 42
rect -599 -30 -593 30
rect -559 -30 -553 30
rect -599 -42 -553 -30
rect -503 30 -457 42
rect -503 -30 -497 30
rect -463 -30 -457 30
rect -503 -42 -457 -30
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect 457 30 503 42
rect 457 -30 463 30
rect 497 -30 503 30
rect 457 -42 503 -30
rect 553 30 599 42
rect 553 -30 559 30
rect 593 -30 599 30
rect 553 -42 599 -30
rect 649 30 695 42
rect 649 -30 655 30
rect 689 -30 695 30
rect 649 -42 695 -30
rect 745 30 791 42
rect 745 -30 751 30
rect 785 -30 791 30
rect 745 -42 791 -30
rect 841 30 887 42
rect 841 -30 847 30
rect 881 -30 887 30
rect 841 -42 887 -30
rect 937 30 983 42
rect 937 -30 943 30
rect 977 -30 983 30
rect 937 -42 983 -30
rect 1033 30 1079 42
rect 1033 -30 1039 30
rect 1073 -30 1079 30
rect 1033 -42 1079 -30
rect 1129 30 1175 42
rect 1129 -30 1135 30
rect 1169 -30 1175 30
rect 1129 -42 1175 -30
rect 1225 30 1271 42
rect 1225 -30 1231 30
rect 1265 -30 1271 30
rect 1225 -42 1271 -30
rect 1321 30 1367 42
rect 1321 -30 1327 30
rect 1361 -30 1367 30
rect 1321 -42 1367 -30
rect 1417 30 1463 42
rect 1417 -30 1423 30
rect 1457 -30 1463 30
rect 1417 -42 1463 -30
rect 1513 30 1559 42
rect 1513 -30 1519 30
rect 1553 -30 1559 30
rect 1513 -42 1559 -30
rect 1609 30 1655 42
rect 1609 -30 1615 30
rect 1649 -30 1655 30
rect 1609 -42 1655 -30
rect 1705 30 1751 42
rect 1705 -30 1711 30
rect 1745 -30 1751 30
rect 1705 -42 1751 -30
rect 1801 30 1847 42
rect 1801 -30 1807 30
rect 1841 -30 1847 30
rect 1801 -42 1847 -30
rect 1897 30 1943 42
rect 1897 -30 1903 30
rect 1937 -30 1943 30
rect 1897 -42 1943 -30
rect 1993 30 2039 42
rect 1993 -30 1999 30
rect 2033 -30 2039 30
rect 1993 -42 2039 -30
rect 2089 30 2135 42
rect 2089 -30 2095 30
rect 2129 -30 2135 30
rect 2089 -42 2135 -30
rect 2185 30 2231 42
rect 2185 -30 2191 30
rect 2225 -30 2231 30
rect 2185 -42 2231 -30
rect 2281 30 2327 42
rect 2281 -30 2287 30
rect 2321 -30 2327 30
rect 2281 -42 2327 -30
rect 2377 30 2423 42
rect 2377 -30 2383 30
rect 2417 -30 2423 30
rect 2377 -42 2423 -30
rect 2473 30 2519 42
rect 2473 -30 2479 30
rect 2513 -30 2519 30
rect 2473 -42 2519 -30
rect 2569 30 2615 42
rect 2569 -30 2575 30
rect 2609 -30 2615 30
rect 2569 -42 2615 -30
rect 2665 30 2711 42
rect 2665 -30 2671 30
rect 2705 -30 2711 30
rect 2665 -42 2711 -30
rect 2761 30 2807 42
rect 2761 -30 2767 30
rect 2801 -30 2807 30
rect 2761 -42 2807 -30
rect 2857 30 2903 42
rect 2857 -30 2863 30
rect 2897 -30 2903 30
rect 2857 -42 2903 -30
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 60 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
