magic
tech sky130A
magscale 1 2
timestamp 1727647182
<< nwell >>
rect -15174 104225 -12341 104240
rect -15174 101448 161454 104225
rect -15174 100934 -12391 101448
rect 2019 101392 161454 101448
rect -15174 -101697 -12341 100934
rect 1348 -9248 1606 -8920
rect 158621 -101697 161454 101392
rect -15174 -104530 161454 -101697
<< pwell >>
rect 1276 -9462 1400 -9306
<< psubdiff >>
rect -18299 107180 -15928 107281
rect 162114 107180 164435 107281
rect -18299 106690 164486 107180
rect -18299 95375 -17534 106690
rect -18198 -102496 -17534 95375
rect -16422 105173 -14905 106690
rect 161678 106286 164486 106690
rect 161678 105173 162589 106286
rect -16422 104758 162589 105173
rect -16422 95375 -15928 104758
rect -16422 -102496 -15964 95375
rect -18198 -104714 -18190 -102496
rect -15972 -104714 -15964 -102496
rect 155796 100790 158000 100809
rect -12010 100168 158000 100790
rect -12010 98854 -11462 100168
rect 155156 99062 158000 100168
rect 155156 98854 156220 99062
rect -12010 98586 156220 98854
rect -11927 97402 -9642 98586
rect -11927 -101312 -11479 97402
rect -10146 -101312 -9642 97402
rect 155796 3296 156220 98586
rect 155768 2849 156220 3296
rect 155768 -2591 156186 2849
rect 155768 -2926 156220 -2591
rect 1308 -9350 1386 -9326
rect 1308 -9424 1332 -9350
rect 1368 -9424 1386 -9350
rect 1308 -9448 1386 -9424
rect 155796 -99116 156220 -2926
rect -11927 -101589 -9642 -101312
rect 17961 -99652 156220 -99116
rect 157553 -98458 158000 99062
rect 157553 -99652 157985 -98458
rect 17961 -99717 157985 -99652
rect 17961 -100983 18676 -99717
rect 46170 -100983 157985 -99717
rect 17961 -101329 157985 -100983
rect 162114 96471 162589 104758
rect -18198 -104916 -17534 -104714
rect -18349 -106504 -17534 -104916
rect -16422 -104916 -15964 -104714
rect 162110 -104916 162589 96471
rect -16422 -105695 162589 -104916
rect -16422 -106504 -15512 -105695
rect -18349 -107212 -15512 -106504
rect 161071 -106908 162589 -105695
rect 163701 104758 164486 106286
rect 163701 94820 164435 104758
rect 163701 -104916 164344 94820
rect 163701 -106908 164486 -104916
rect 161071 -107212 164486 -106908
rect -18349 -107893 164486 -107212
<< nsubdiff >>
rect -14661 103067 158938 103707
rect -14661 102035 -14169 103067
rect 158791 102035 158938 103067
rect -14661 101691 158938 102035
rect 159086 102674 161151 103903
rect -14611 101101 -12743 101691
rect -14611 95717 -14316 101101
rect -14735 92859 -14316 95717
rect -14611 -101810 -14316 92859
rect -14647 -103373 -14316 -101810
rect -13136 -101810 -12743 101101
rect 1394 -8986 1554 -8958
rect 1394 -9176 1440 -8986
rect 1518 -9176 1554 -8986
rect 1394 -9206 1554 -9176
rect 159086 -101702 159578 102674
rect 160659 -101702 161151 102674
rect 159086 -101810 161151 -101702
rect -13136 -102411 161151 -101810
rect -13136 -103373 -11982 -102411
rect -14647 -103513 -11982 -103373
rect 159874 -103513 161151 -102411
rect -14647 -104003 161151 -103513
rect 159086 -104013 161151 -104003
<< psubdiffcont >>
rect -17534 -102496 -16422 106690
rect -14905 105173 161678 106690
rect -18190 -104714 -15972 -102496
rect -11462 98854 155156 100168
rect -11479 -101312 -10146 97402
rect 156220 2849 157553 99062
rect 156186 -2591 157553 2849
rect 1332 -9424 1368 -9350
rect 156220 -99652 157553 -2591
rect 18676 -100983 46170 -99717
rect -17534 -106504 -16422 -104714
rect -15512 -107212 161071 -105695
rect 162589 -106908 163701 106286
<< nsubdiffcont >>
rect -14169 102035 158791 103067
rect -14316 -103373 -13136 101101
rect 1440 -9176 1518 -8986
rect 159578 -101702 160659 102674
rect -11982 -103513 159874 -102411
<< poly >>
rect 14511 3294 14739 3313
rect 14511 3230 14534 3294
rect 14608 3285 14739 3294
rect 14608 3231 15303 3285
rect 14608 3230 14739 3231
rect 14511 3217 14739 3230
rect 148146 1776 148244 1796
rect 148146 1456 148162 1776
rect 148228 1456 148244 1776
rect 148146 1248 148244 1456
rect 148148 562 148246 1124
rect 148150 238 148248 344
rect 148150 136 148170 238
rect 148230 136 148248 238
rect 148150 110 148248 136
rect 14428 -3836 14539 -3806
rect 14428 -3904 14451 -3836
rect 14509 -3837 14539 -3836
rect 14602 -3837 15223 -3836
rect 14509 -3893 15223 -3837
rect 14509 -3895 14634 -3893
rect 14509 -3904 14539 -3895
rect 14428 -3927 14539 -3904
<< polycont >>
rect 14534 3230 14608 3294
rect 148162 1456 148228 1776
rect 148170 136 148230 238
rect 14451 -3904 14509 -3836
<< locali >>
rect -18299 107180 -15928 107281
rect 162114 107180 164435 107281
rect -18299 106690 164486 107180
rect -18299 95375 -17534 106690
rect -22430 3452 -18535 3469
rect -22430 3207 -18510 3452
rect -22430 2324 -22119 3207
rect -19207 2324 -18510 3207
rect -22430 2075 -18510 2324
rect -18918 -110654 -18510 2075
rect -18198 -102496 -17534 95375
rect -18198 -104714 -18190 -102496
rect -18198 -104916 -17534 -104714
rect -18349 -106504 -17534 -104916
rect -16422 105173 -14905 106690
rect 161678 106286 164486 106690
rect 161678 105173 162589 106286
rect -16422 104758 162589 105173
rect -16422 95375 -15928 104758
rect -14736 103067 160953 103736
rect -14736 102035 -14169 103067
rect 158791 102772 160953 103067
rect 158791 102035 159528 102772
rect -14736 101866 159528 102035
rect -14736 101101 -12705 101866
rect -16422 -102496 -15964 95375
rect -14736 94984 -14316 101101
rect -14735 92859 -14316 94984
rect -15972 -104714 -15964 -102496
rect -14575 -103373 -14316 92859
rect -13136 -102107 -12705 101101
rect -11927 100718 -9642 100756
rect -11927 100168 158008 100718
rect -11927 98854 -11462 100168
rect 155156 99062 158008 100168
rect 155156 98854 156220 99062
rect -11927 98538 156220 98854
rect -11927 97402 -9642 98538
rect -11927 -101312 -11479 97402
rect -10146 -101312 -9642 97402
rect 14511 3294 14633 3313
rect 155793 3296 156220 98538
rect 14511 3230 14534 3294
rect 14608 3230 14633 3294
rect 14511 3217 14633 3230
rect 155768 2849 156220 3296
rect 157553 98538 158008 99062
rect 148148 1776 148248 1794
rect 148148 1456 148162 1776
rect 148228 1456 148248 1776
rect 148148 1440 148248 1456
rect 148150 238 148244 254
rect 148150 136 148170 238
rect 148230 136 148244 238
rect 148150 110 148244 136
rect 155768 -2591 156186 2849
rect 155768 -2926 156220 -2591
rect 14428 -3836 14539 -3806
rect 14428 -3904 14451 -3836
rect 14509 -3904 14539 -3836
rect 14428 -3927 14539 -3904
rect 1244 -8980 1556 -8944
rect 1394 -8986 1554 -8980
rect 1394 -9176 1440 -8986
rect 1518 -9176 1554 -8986
rect 1394 -9206 1554 -9176
rect 1258 -9246 1368 -9244
rect 1194 -9250 1368 -9246
rect 626 -9276 992 -9260
rect 626 -9336 646 -9276
rect 962 -9285 992 -9276
rect 962 -9331 1158 -9285
rect 1194 -9286 1274 -9250
rect 1352 -9286 1368 -9250
rect 1194 -9292 1368 -9286
rect 962 -9336 992 -9331
rect 626 -9350 992 -9336
rect 1308 -9350 1386 -9326
rect 1308 -9424 1332 -9350
rect 1368 -9424 1386 -9350
rect 1308 -9434 1386 -9424
rect 1224 -9444 1386 -9434
rect 1218 -9482 1386 -9444
rect 1218 -9492 1380 -9482
rect 155793 -99106 156220 -2926
rect 44154 -99133 156220 -99106
rect -11927 -101589 -9642 -101312
rect 17972 -99652 156220 -99133
rect 157553 -99106 157979 98538
rect 157553 -99652 157983 -99106
rect 17972 -99698 157983 -99652
rect 17972 -99717 42624 -99698
rect 17972 -99736 18676 -99717
rect 17972 -100999 18658 -99736
rect 157466 -100999 157983 -99698
rect 17972 -101356 157983 -100999
rect 155793 -101388 157979 -101356
rect 159083 -101702 159528 101866
rect 160708 -101702 160953 102772
rect 162114 96471 162589 104758
rect 159083 -102107 160953 -101702
rect -13136 -102411 160953 -102107
rect -13136 -103373 -11982 -102411
rect -14575 -103513 -11982 -103373
rect 159874 -103513 160953 -102411
rect -14575 -103977 160953 -103513
rect -16422 -104916 -15964 -104714
rect 162110 -104916 162589 96471
rect -16422 -105695 162589 -104916
rect -16422 -106504 -15512 -105695
rect -18349 -107212 -15512 -106504
rect 161071 -106908 162589 -105695
rect 163701 104758 164486 106286
rect 163701 94820 164435 104758
rect 163701 -104916 164344 94820
rect 163701 -106908 164486 -104916
rect 161071 -107212 164486 -106908
rect -18349 -107893 164486 -107212
rect -18918 -110928 -12069 -110654
rect -18918 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18918 -111995 -12069 -111747
rect -18918 -112075 -18510 -111995
<< viali >>
rect -22119 2324 -19207 3207
rect -17534 -106504 -16422 106690
rect -14905 105173 161678 106690
rect -14169 102035 158791 103067
rect 159528 102674 160708 102772
rect -14316 -103373 -13136 101101
rect -11462 98854 155156 100168
rect -11479 -101312 -10146 97402
rect 14534 3230 14608 3294
rect 156220 2849 157553 99062
rect 148162 1456 148228 1776
rect 148170 136 148230 238
rect 156186 -2591 157553 2849
rect 14451 -3904 14509 -3836
rect 646 -9336 962 -9276
rect 1274 -9286 1352 -9250
rect 156220 -99652 157553 -2591
rect 42624 -99717 157466 -99698
rect 42624 -99736 46170 -99717
rect 18658 -100983 18676 -99736
rect 18676 -100983 46170 -99736
rect 46170 -100983 157466 -99717
rect 18658 -100999 157466 -100983
rect 159528 -101702 159578 102674
rect 159578 -101702 160659 102674
rect 160659 -101702 160708 102674
rect -11982 -103513 159874 -102411
rect -15512 -107212 161071 -105695
rect 162589 -106908 163701 106286
rect -18327 -111747 -12516 -110928
<< metal1 >>
rect -18299 107180 -15928 107281
rect 162114 107180 164435 107281
rect -18299 106690 164486 107180
rect -18299 95375 -17534 106690
rect -22408 3207 -18497 3481
rect -22408 2324 -22119 3207
rect -19207 2324 -18497 3207
rect -22408 2088 -18497 2324
rect -18198 -104916 -17534 95375
rect -18349 -106504 -17534 -104916
rect -16422 105173 -14905 106690
rect 161678 106286 164486 106690
rect 161678 105173 162589 106286
rect -16422 104758 162589 105173
rect -16422 95375 -15928 104758
rect -14653 103671 161041 103760
rect -14653 103067 161066 103671
rect -14653 102035 -14169 103067
rect 158791 102772 161066 103067
rect 158791 102035 159528 102772
rect -14653 101808 159528 102035
rect -14646 101101 -12798 101808
rect -14646 96938 -14316 101101
rect -14725 95717 -14316 96938
rect -16422 -104916 -15964 95375
rect -14735 92859 -14316 95717
rect -14646 -103373 -14316 92859
rect -13136 96938 -12798 101101
rect -11927 100718 -9642 100756
rect -11927 100168 158008 100718
rect -11927 98854 -11462 100168
rect 155156 99062 158008 100168
rect 155156 98854 156220 99062
rect -11927 98538 156220 98854
rect -11927 97402 -9642 98538
rect -13136 92863 -12747 96938
rect -13136 -102046 -12798 92863
rect -11927 -101312 -11479 97402
rect -10146 -99709 -9642 97402
rect -42 48182 794 48218
rect -42 48122 62 48182
rect 736 48122 794 48182
rect -42 48072 794 48122
rect -3767 48070 794 48072
rect -6574 47862 794 48070
rect -6574 46716 -3222 47862
rect -42 47860 794 47862
rect -3782 -2028 -3222 46716
rect -3782 -5352 -3614 -2028
rect -3246 -5352 -3222 -2028
rect -3782 -48482 -3222 -5352
rect -3052 46322 -2492 46326
rect -3052 46280 800 46322
rect -3052 46222 44 46280
rect 766 46222 800 46280
rect -3052 46180 800 46222
rect -3052 -6518 -2492 46180
rect -2380 44396 -1820 44402
rect 0 44396 800 44412
rect -2380 44386 800 44396
rect -2380 44368 28 44386
rect -2380 44230 -1820 44368
rect 0 44328 28 44368
rect 746 44328 800 44386
rect 0 44298 800 44328
rect -2380 42908 -2286 44230
rect -1922 42908 -1820 44230
rect -2380 37720 -1820 42908
rect -1693 42494 -1142 42502
rect -12 42494 816 42502
rect -1694 42476 816 42494
rect -1694 42418 78 42476
rect 742 42418 816 42476
rect -1694 42390 816 42418
rect -1694 42376 810 42390
rect -1693 41992 -1142 42376
rect -1693 41586 -1588 41992
rect -1702 40534 -1588 41586
rect -1224 40534 -1142 41992
rect -2380 37692 -1982 37720
rect -3052 -7226 -2964 -6518
rect -2554 -7226 -2492 -6518
rect -3052 -7300 -2492 -7226
rect -2380 35774 -1964 35776
rect -2380 35554 -1820 35774
rect -2380 33956 -2262 35554
rect -1926 33956 -1820 35554
rect -3052 -8660 -2492 -8508
rect -3052 -9368 -2964 -8660
rect -2554 -9368 -2492 -8660
rect -3052 -46794 -2492 -9368
rect -2380 -44988 -1820 33956
rect -1702 -43000 -1142 40534
rect -1034 40608 -474 40610
rect -1034 40566 794 40608
rect -1034 40510 64 40566
rect 738 40510 794 40566
rect -1034 40456 794 40510
rect -1034 39544 -474 40456
rect -1034 38202 -1026 39544
rect -526 38202 -474 39544
rect -352 38708 208 38712
rect -354 38664 794 38708
rect -354 38598 66 38664
rect 716 38598 794 38664
rect -354 38572 794 38598
rect -1034 -41096 -474 38202
rect -352 -8140 208 38572
rect 8660 4060 9130 4316
rect 10226 4194 10552 4358
rect 3294 3212 4770 3444
rect 8660 3350 8916 4060
rect 3294 2288 3492 3212
rect 4532 2288 4770 3212
rect 8606 3276 8962 3350
rect 8606 2824 8662 3276
rect 8896 2824 8962 3276
rect 8606 2784 8962 2824
rect 8730 2782 8802 2784
rect 9942 2638 10100 2996
rect 3294 2068 4770 2288
rect 9938 2606 10100 2638
rect 786 1027 948 1055
rect 786 912 811 1027
rect 922 980 948 1027
rect 922 978 2505 980
rect 922 966 2534 978
rect 922 938 2394 966
rect 922 912 948 938
rect 786 887 948 912
rect 1092 912 2394 938
rect 2504 912 2534 966
rect 1092 896 2534 912
rect 3878 -270 4023 2068
rect 9938 730 10038 2606
rect 10388 2256 10552 4194
rect 12492 4212 13874 4296
rect 12492 3792 12636 4212
rect 13752 3792 13874 4212
rect 12492 3768 13874 3792
rect 148142 3818 148242 3900
rect 12492 3714 14926 3768
rect 13344 3706 14926 3714
rect 148142 3732 151160 3818
rect 14374 2792 14482 3537
rect 148142 3528 148252 3732
rect 151036 3528 151160 3732
rect 148142 3436 151160 3528
rect 14511 3294 14633 3313
rect 14511 3230 14534 3294
rect 14608 3230 14633 3294
rect 14511 3217 14633 3230
rect 14870 3274 15020 3292
rect 14870 3222 14923 3274
rect 15006 3262 15020 3274
rect 15006 3222 15086 3262
rect 14870 3206 15086 3222
rect 14870 3205 15020 3206
rect 14983 2912 15595 2991
rect 14236 2774 14682 2792
rect 14236 2720 14683 2774
rect 14236 2396 14298 2720
rect 14596 2710 14683 2720
rect 14596 2396 14682 2710
rect 14983 2678 15073 2912
rect 15496 2678 15595 2912
rect 14983 2604 15595 2678
rect 14236 2318 14682 2396
rect 10346 2186 10626 2256
rect 10346 1902 10408 2186
rect 10572 1902 10626 2186
rect 10346 1848 10626 1902
rect 148142 1798 148242 3436
rect 155793 3296 156220 98538
rect 155768 2849 156220 3296
rect 157553 98538 158008 99062
rect 151204 1946 152196 2020
rect 148142 1776 148244 1798
rect 148142 1456 148162 1776
rect 148228 1456 148244 1776
rect 151204 1770 151268 1946
rect 152032 1770 152196 1946
rect 151204 1725 152196 1770
rect 151208 1574 151548 1725
rect 151674 1567 152013 1725
rect 148142 1438 148244 1456
rect 141714 868 143268 950
rect 148100 945 148136 1242
rect 148264 1160 148394 1168
rect 148264 1138 148320 1160
rect 148254 1108 148320 1138
rect 148384 1108 148394 1160
rect 148254 1104 148394 1108
rect 148264 1098 148394 1104
rect 148264 1096 148346 1098
rect 9932 698 10060 730
rect 7468 630 8208 670
rect 7554 582 7658 602
rect 7554 274 7582 582
rect 7358 260 7582 274
rect 7642 260 7658 582
rect 7358 234 7658 260
rect 7358 232 7634 234
rect 4212 -106 4364 -90
rect 4212 -168 4242 -106
rect 4326 -168 4364 -106
rect 4212 -178 4364 -168
rect 3878 -304 4136 -270
rect 3974 -314 4136 -304
rect 3974 -316 4023 -314
rect 6970 -428 7064 -94
rect 6820 -472 7064 -428
rect 6820 -556 6880 -472
rect 7024 -556 7064 -472
rect 6820 -606 7064 -556
rect 5690 -782 5782 -764
rect 5088 -852 5250 -844
rect 5088 -904 5110 -852
rect 5216 -862 5250 -852
rect 5216 -904 5428 -862
rect 5088 -910 5428 -904
rect 5690 -894 5708 -782
rect 5768 -894 5782 -782
rect 5690 -910 5782 -894
rect 5088 -916 5250 -910
rect 8064 -4072 8208 630
rect 9932 562 9956 698
rect 10042 562 10060 698
rect 9932 536 10060 562
rect 9938 462 10038 536
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 147518 905 148136 945
rect 147518 791 147540 905
rect 147666 791 148136 905
rect 147518 754 148136 791
rect 141714 440 143268 508
rect 148100 496 148136 754
rect 10076 -66 10462 40
rect 10076 -380 10164 -66
rect 10374 -236 10462 -66
rect 141923 -176 142237 440
rect 148259 384 148298 543
rect 148257 345 148437 384
rect 148150 238 148244 254
rect 148150 136 148170 238
rect 148230 136 148244 238
rect 148150 110 148244 136
rect 10374 -242 14172 -236
rect 10374 -264 14792 -242
rect 10374 -380 14078 -264
rect 10076 -382 14078 -380
rect 14758 -382 14792 -264
rect 10076 -394 14792 -382
rect 10076 -402 14172 -394
rect 10076 -526 10462 -402
rect 15072 -490 147551 -176
rect 148398 -2319 148437 345
rect 151372 382 151468 388
rect 151372 308 151384 382
rect 151456 308 151468 382
rect 151372 296 151468 308
rect 153290 366 153432 394
rect 150720 174 151114 214
rect 150720 68 150748 174
rect 151082 68 151114 174
rect 150720 46 151114 68
rect 151950 -83 152126 -74
rect 151950 -90 152127 -83
rect 151950 -158 151964 -90
rect 152116 -158 152127 -90
rect 151950 -170 152127 -158
rect 152073 -690 152127 -170
rect 152790 -782 152940 192
rect 153290 120 153310 366
rect 153414 120 153432 366
rect 153290 100 153432 120
rect 148384 -2336 154888 -2319
rect 148384 -2375 154901 -2336
rect 148384 -2535 154888 -2375
rect 148384 -2736 154896 -2535
rect 148400 -2952 154896 -2736
rect 155768 -2591 156186 2849
rect 155768 -2926 156220 -2591
rect 14666 -3198 15268 -3130
rect 10457 -3600 10626 -3454
rect 10894 -3493 14103 -3454
rect 10456 -3618 10854 -3600
rect 10894 -3618 14007 -3493
rect 10456 -3666 14007 -3618
rect 10456 -3898 10526 -3666
rect 10794 -3742 14007 -3666
rect 14068 -3742 14103 -3493
rect 14666 -3504 14748 -3198
rect 15165 -3504 15268 -3198
rect 14666 -3599 15268 -3504
rect 10794 -3764 14103 -3742
rect 10794 -3898 10854 -3764
rect 14799 -3800 15016 -3768
rect 10456 -3966 10854 -3898
rect 14428 -3836 14539 -3806
rect 14428 -3904 14451 -3836
rect 14509 -3904 14539 -3836
rect 14428 -3927 14539 -3904
rect 14799 -3906 14836 -3800
rect 14948 -3815 15016 -3800
rect 14948 -3849 15346 -3815
rect 14948 -3906 15016 -3849
rect 14799 -3935 15016 -3906
rect 7680 -4148 8400 -4072
rect 7680 -4390 7776 -4148
rect 8296 -4390 8400 -4148
rect 7680 -4456 8400 -4390
rect 10457 -6322 10767 -3966
rect 12980 -4086 13876 -3948
rect 12980 -4494 13094 -4086
rect 13714 -4314 13876 -4086
rect 14543 -4187 14579 -4077
rect 15400 -4187 16157 -4186
rect 14543 -4223 14586 -4187
rect 15358 -4223 16157 -4187
rect 13714 -4392 13893 -4314
rect 13714 -4494 13876 -4392
rect 12980 -4572 13876 -4494
rect 14543 -4666 14579 -4223
rect 15400 -4227 16157 -4223
rect 15400 -4348 15558 -4227
rect 15997 -4348 16157 -4227
rect 15400 -4387 16157 -4348
rect 14300 -4744 14624 -4666
rect 14300 -4954 14392 -4744
rect 14550 -4954 14624 -4744
rect 14300 -5036 14624 -4954
rect 10994 -5486 11342 -5446
rect 10994 -5800 11040 -5486
rect 11300 -5800 11342 -5486
rect 10994 -5834 11342 -5800
rect 10458 -6498 10767 -6322
rect 10474 -6508 10767 -6498
rect 11057 -7643 11091 -5834
rect 11057 -7677 11528 -7643
rect -352 -8190 783 -8140
rect -352 -39194 208 -8190
rect 2658 -8472 2742 -8464
rect 2656 -8532 2742 -8472
rect 1284 -8978 1664 -8914
rect 1284 -9042 1330 -8978
rect 1618 -9042 1664 -8978
rect 1284 -9066 1664 -9042
rect 2656 -9108 2820 -8532
rect 2234 -9144 2820 -9108
rect 9222 -9122 9272 -8930
rect 11486 -9122 11558 -8901
rect 1812 -9236 1938 -9228
rect 1258 -9246 1368 -9244
rect 1812 -9246 1832 -9236
rect 1196 -9250 1832 -9246
rect 626 -9276 992 -9260
rect 626 -9336 646 -9276
rect 962 -9336 992 -9276
rect 1196 -9286 1274 -9250
rect 1352 -9286 1832 -9250
rect 1196 -9290 1832 -9286
rect 1920 -9290 1938 -9236
rect 1196 -9292 1938 -9290
rect 1812 -9294 1938 -9292
rect 626 -9350 992 -9336
rect 1650 -9494 1976 -9424
rect 2234 -9494 2270 -9144
rect 2656 -9158 2820 -9144
rect 2656 -9194 3014 -9158
rect 8594 -9194 11558 -9122
rect 1212 -9530 2270 -9494
rect 1650 -9617 1976 -9530
rect 497 -9682 1976 -9617
rect 497 -9892 526 -9682
rect 1804 -9892 1976 -9682
rect 497 -9943 1976 -9892
rect -352 -39220 472 -39194
rect -352 -39290 -276 -39220
rect 422 -39290 472 -39220
rect -352 -39314 472 -39290
rect -352 -39336 208 -39314
rect -1036 -41120 476 -41096
rect -1036 -41188 -260 -41120
rect 424 -41188 476 -41120
rect -1036 -41216 476 -41188
rect -1034 -41224 -474 -41216
rect -1704 -43030 472 -43000
rect -1704 -43088 -262 -43030
rect 436 -43088 472 -43030
rect -1704 -43124 472 -43088
rect -1702 -43128 -1142 -43124
rect -314 -44940 472 -44906
rect -314 -44988 -284 -44940
rect -2380 -45004 -284 -44988
rect 436 -45004 472 -44940
rect -2380 -45006 472 -45004
rect -2360 -45016 472 -45006
rect -314 -45032 472 -45016
rect -3052 -46846 474 -46794
rect -3052 -46904 -248 -46846
rect 416 -46904 474 -46846
rect -3052 -46936 474 -46904
rect -3052 -46956 -2492 -46936
rect -3782 -48692 545 -48482
rect -336 -48748 542 -48692
rect -336 -48810 -298 -48748
rect 442 -48810 542 -48748
rect -336 -48836 542 -48810
rect 155793 -99080 156220 -2926
rect 10473 -99429 14022 -99129
rect 10473 -99709 10773 -99429
rect -10146 -100779 10773 -99709
rect 13547 -99754 14022 -99429
rect 17949 -99652 156220 -99080
rect 157553 -99120 157979 98538
rect 157553 -99652 157985 -99120
rect 17949 -99698 157985 -99652
rect 17949 -99709 42624 -99698
rect 15947 -99736 42624 -99709
rect 15947 -99754 18658 -99736
rect 13547 -100779 18658 -99754
rect -10146 -100999 18658 -100779
rect 157466 -100999 157985 -99698
rect -10146 -101081 157985 -100999
rect -10146 -101312 -9642 -101081
rect 9573 -101104 17446 -101081
rect -11927 -101589 -9642 -101312
rect 17949 -101360 157985 -101081
rect 17949 -101379 157979 -101360
rect 155793 -101388 157979 -101379
rect 159224 -101702 159528 101808
rect 160708 -101702 161066 102772
rect 162114 96471 162589 104758
rect 159224 -102046 161066 -101702
rect -13136 -102104 10523 -102046
rect 15947 -102104 161066 -102046
rect -13136 -102411 161066 -102104
rect -13136 -103373 -11982 -102411
rect -14646 -103513 -11982 -103373
rect 159874 -103513 161066 -102411
rect -14646 -103958 161066 -103513
rect -14513 -103963 161066 -103958
rect 159224 -103989 161066 -103963
rect 162110 -104916 162589 96471
rect -16422 -105681 162589 -104916
rect -16422 -105695 10989 -105681
rect 13851 -105695 162589 -105681
rect -16422 -106504 -15512 -105695
rect -18349 -107212 -15512 -106504
rect 161071 -106908 162589 -105695
rect 163701 104758 164486 106286
rect 163701 94820 164435 104758
rect 163701 -104916 164344 94820
rect 163701 -106908 164486 -104916
rect 161071 -107212 164486 -106908
rect -18349 -107252 10989 -107212
rect 13851 -107252 164486 -107212
rect -18349 -107893 164486 -107252
rect -18198 -108095 -15964 -107893
rect -18798 -110928 -12069 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18798 -111995 -12069 -111747
<< via1 >>
rect -22119 2324 -19207 3207
rect 62 48122 736 48182
rect -3614 -5352 -3246 -2028
rect 44 46222 766 46280
rect 28 44328 746 44386
rect -2286 42908 -1922 44230
rect 78 42418 742 42476
rect -1588 40534 -1224 41992
rect -2964 -7226 -2554 -6518
rect -2262 33956 -1926 35554
rect -2964 -9368 -2554 -8660
rect 64 40510 738 40566
rect -1026 38202 -526 39544
rect 66 38598 716 38664
rect 3492 2288 4532 3212
rect 8662 2824 8896 3276
rect 811 912 922 1027
rect 2394 912 2504 966
rect 12636 3792 13752 4212
rect 148252 3528 151036 3732
rect 14534 3230 14608 3294
rect 14923 3222 15006 3274
rect 14298 2396 14596 2720
rect 15073 2678 15496 2912
rect 10408 1902 10572 2186
rect 151268 1770 152032 1946
rect 148320 1108 148384 1160
rect 7582 260 7642 582
rect 4242 -168 4326 -106
rect 6880 -556 7024 -472
rect 5110 -904 5216 -852
rect 5708 -894 5768 -782
rect 9956 562 10042 698
rect 141758 508 143186 868
rect 147540 791 147666 905
rect 10164 -380 10374 -66
rect 148170 136 148230 238
rect 14078 -382 14758 -264
rect 151384 308 151456 382
rect 150748 68 151082 174
rect 151964 -158 152116 -90
rect 153310 120 153414 366
rect 10526 -3898 10794 -3666
rect 14007 -3742 14068 -3493
rect 14748 -3504 15165 -3198
rect 14451 -3904 14509 -3836
rect 14836 -3906 14948 -3800
rect 7776 -4390 8296 -4148
rect 13094 -4494 13714 -4086
rect 15558 -4348 15997 -4227
rect 14392 -4954 14550 -4744
rect 11040 -5800 11300 -5486
rect 1330 -9042 1618 -8978
rect 646 -9336 962 -9276
rect 1832 -9290 1920 -9236
rect 526 -9892 1804 -9682
rect -276 -39290 422 -39220
rect -260 -41188 424 -41120
rect -262 -43088 436 -43030
rect -284 -45004 436 -44940
rect -248 -46904 416 -46846
rect -298 -48810 442 -48748
rect 10773 -100779 13547 -99429
rect 159607 1871 160669 3056
rect 10989 -105695 13851 -105681
rect 10989 -107212 13851 -105695
rect 10989 -107252 13851 -107212
rect -18327 -111747 -12516 -110928
<< metal2 >>
rect 133308 87497 148018 87509
rect 133308 87428 148020 87497
rect 133308 87269 166338 87428
rect 146558 79019 166338 87269
rect -2 48182 794 48220
rect -2 48122 62 48182
rect 736 48122 794 48182
rect -2 48094 794 48122
rect -2 46280 802 46310
rect -2 46222 44 46280
rect 766 46222 802 46280
rect -2 46192 802 46222
rect 0 44386 800 44412
rect -8551 44230 -1816 44386
rect 0 44328 28 44386
rect 746 44328 800 44386
rect 0 44298 800 44328
rect -8551 42908 -2286 44230
rect -1922 42908 -1816 44230
rect -8551 42824 -1816 42908
rect -12 42476 816 42502
rect -12 42418 78 42476
rect 742 42418 816 42476
rect -12 42390 816 42418
rect -8468 41992 -1150 42074
rect -8468 40534 -1588 41992
rect -1224 40534 -1150 41992
rect -8468 40388 -1150 40534
rect 2 40566 788 40606
rect 2 40510 64 40566
rect 738 40510 788 40566
rect 2 40484 788 40510
rect -8260 39544 -494 39628
rect -8260 38202 -1026 39544
rect -526 38202 -494 39544
rect 0 38664 784 38692
rect 0 38598 66 38664
rect 716 38598 784 38664
rect 0 38576 784 38598
rect -8260 38108 -494 38202
rect -2372 35554 -1814 35752
rect -2372 33956 -2262 35554
rect -1926 33956 -1814 35554
rect -2372 33750 -1814 33956
rect -4264 4744 890 7690
rect 8568 6950 11198 7294
rect 7701 6536 7742 6772
rect 8568 6536 8960 6950
rect 7701 6530 8960 6536
rect 7684 6495 8960 6530
rect -22408 3207 -18497 3481
rect -22408 2324 -22119 3207
rect -19207 2324 -18497 3207
rect -22408 2088 -18497 2324
rect -2626 3266 -1628 4744
rect -2626 2398 -2468 3266
rect -1848 2398 -1628 3266
rect -2626 2132 -1628 2398
rect 3294 3212 4770 3444
rect 3294 2288 3492 3212
rect 4532 2288 4770 3212
rect 3294 2068 4770 2288
rect -5184 -680 674 1248
rect 786 1027 948 1055
rect 786 912 811 1027
rect 922 912 948 1027
rect 2381 982 2459 985
rect 786 887 948 912
rect 2374 966 2524 982
rect 2374 912 2394 966
rect 2504 912 2524 966
rect 2374 -94 2524 912
rect 7684 636 7864 6495
rect 8568 5410 8960 6495
rect 10878 5410 11198 6950
rect 8568 5070 11198 5410
rect 10674 4572 11058 5070
rect 10677 4130 11058 4572
rect 10674 3980 11058 4130
rect 8606 3276 8962 3350
rect 8606 2824 8662 3276
rect 8896 2824 8962 3276
rect 8606 2784 8962 2824
rect 10668 3172 11058 3980
rect 12520 4212 13874 4286
rect 12520 3792 12636 4212
rect 13752 3792 13874 4212
rect 12520 3712 13874 3792
rect 148146 3732 151160 3818
rect 148146 3528 148252 3732
rect 151036 3528 151160 3732
rect 148146 3436 151160 3528
rect 14052 3294 14634 3313
rect 14051 3230 14534 3294
rect 14608 3230 14634 3294
rect 14051 3217 14634 3230
rect 14870 3274 15020 3292
rect 14870 3222 14923 3274
rect 15006 3262 15020 3274
rect 15833 3272 16533 3315
rect 15006 3261 15086 3262
rect 15833 3261 15888 3272
rect 15006 3222 15888 3261
rect 14051 3172 14162 3217
rect 14870 3206 15888 3222
rect 14870 3205 15020 3206
rect 15833 3184 15888 3206
rect 16384 3184 16533 3272
rect 10668 2940 14163 3172
rect 15833 3149 16533 3184
rect 159058 3056 161125 3278
rect 10346 2186 10626 2256
rect 10346 1902 10408 2186
rect 10572 1902 10626 2186
rect 10346 1848 10626 1902
rect 10668 1512 11058 2940
rect 14983 2912 15595 2991
rect 148400 2983 148817 3023
rect 14236 2735 14374 2792
rect 14482 2735 14682 2792
rect 14236 2720 14682 2735
rect 14236 2396 14298 2720
rect 14596 2396 14682 2720
rect 14983 2678 15073 2912
rect 15496 2678 15595 2912
rect 14983 2604 15595 2678
rect 148370 2667 154640 2983
rect 148370 2566 154648 2667
rect 14236 2318 14682 2396
rect 148378 2250 154648 2566
rect 7554 582 7658 602
rect 7554 260 7582 582
rect 7642 260 7658 582
rect 7554 234 7658 260
rect 7560 232 7634 234
rect 7694 204 7864 636
rect 9932 698 10060 730
rect 9932 562 9956 698
rect 10042 562 10060 698
rect 9932 536 10060 562
rect 2374 -106 4362 -94
rect 2374 -168 4242 -106
rect 4326 -168 4362 -106
rect 2374 -172 4362 -168
rect 6820 -472 7064 -428
rect 6820 -556 6880 -472
rect 7024 -556 7064 -472
rect 6820 -606 7064 -556
rect -5108 -906 -4096 -680
rect 5690 -782 5782 -764
rect -5108 -1554 -4990 -906
rect -4196 -1554 -4096 -906
rect 4570 -848 4732 -832
rect 4570 -916 4588 -848
rect 4714 -862 4732 -848
rect 5088 -852 5250 -844
rect 5088 -862 5110 -852
rect 4714 -904 5110 -862
rect 5216 -904 5250 -852
rect 4714 -912 5250 -904
rect 5690 -894 5708 -782
rect 5768 -894 5782 -782
rect 5690 -910 5782 -894
rect 4714 -916 4732 -912
rect 5088 -916 5250 -912
rect 4570 -932 4732 -916
rect 7684 -1294 7864 204
rect 10076 -66 10462 40
rect 10076 -380 10164 -66
rect 10374 -380 10462 -66
rect 10076 -526 10462 -380
rect 10668 -806 11056 1512
rect 148383 1168 148425 2250
rect 151204 2019 152196 2020
rect 159058 2019 159607 3056
rect 151203 1946 159607 2019
rect 151203 1770 151268 1946
rect 152032 1871 159607 1946
rect 160669 2019 161125 3056
rect 160669 1871 161171 2019
rect 152032 1770 161171 1871
rect 151203 1680 161171 1770
rect 148312 1160 148425 1168
rect 148312 1138 148320 1160
rect 148254 1108 148320 1138
rect 148384 1108 148425 1160
rect 148254 1104 148425 1108
rect 148312 1098 148425 1104
rect 148383 1097 148425 1098
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 147518 905 147705 945
rect 147518 791 147540 905
rect 147666 791 147705 905
rect 147518 754 147705 791
rect 141714 440 143268 508
rect 142442 156 142662 440
rect 151372 382 151468 390
rect 151372 308 151384 382
rect 151456 308 151468 382
rect 148148 238 148244 304
rect 12778 -64 147436 156
rect 148148 136 148170 238
rect 148230 142 148244 238
rect 150720 174 151114 214
rect 148230 136 148414 142
rect 148148 46 148414 136
rect 150720 68 150748 174
rect 151082 68 151114 174
rect 150720 46 151114 68
rect 151372 -74 151468 308
rect 153288 366 153436 396
rect 153288 120 153310 366
rect 153414 120 153436 366
rect 151372 -90 152128 -74
rect 151372 -158 151964 -90
rect 152116 -158 152128 -90
rect 151372 -170 152128 -158
rect 14046 -244 14792 -242
rect 153288 -244 153436 120
rect 14046 -264 153436 -244
rect 14046 -382 14078 -264
rect 14758 -382 153436 -264
rect 14046 -392 153436 -382
rect 14046 -394 14792 -392
rect 10088 -894 11056 -806
rect 12788 -808 150818 -588
rect -5108 -1672 -4096 -1554
rect -3754 -2028 -3176 -1728
rect -3754 -4654 -3614 -2028
rect -3766 -4766 -3614 -4654
rect -3778 -4966 -3614 -4766
rect -3754 -5352 -3614 -4966
rect -3246 -4654 -3176 -2028
rect 8528 -2976 9800 -2932
rect 8528 -3338 8576 -2976
rect 9764 -3338 9800 -2976
rect 8528 -3380 9800 -3338
rect 7680 -4148 8400 -4072
rect 7680 -4390 7776 -4148
rect 8296 -4390 8400 -4148
rect 7680 -4456 8400 -4390
rect -3246 -4712 9218 -4654
rect -3246 -4916 8224 -4712
rect 9050 -4916 9218 -4712
rect -3246 -4966 9218 -4916
rect -3246 -5352 -3176 -4966
rect -3754 -5514 -3176 -5352
rect 10091 -6056 10344 -894
rect 150598 -1836 150818 -808
rect 152818 -1836 153038 -1276
rect 150598 -2056 153038 -1836
rect 14666 -3198 15268 -3130
rect 13967 -3493 14098 -3453
rect 10456 -3666 10854 -3600
rect 10456 -3898 10526 -3666
rect 10794 -3898 10854 -3666
rect 10456 -3966 10854 -3898
rect 13967 -3742 14007 -3493
rect 14068 -3742 14098 -3493
rect 14666 -3504 14748 -3198
rect 15165 -3504 15268 -3198
rect 14666 -3599 15268 -3504
rect 13967 -3806 14098 -3742
rect 14799 -3800 16230 -3769
rect 13967 -3836 14539 -3806
rect 13967 -3904 14451 -3836
rect 14509 -3904 14539 -3836
rect 13967 -3927 14539 -3904
rect 14799 -3906 14836 -3800
rect 14948 -3906 16230 -3800
rect 13967 -3929 14520 -3927
rect 13967 -3932 14202 -3929
rect 14799 -3935 16230 -3906
rect 12980 -4086 13876 -3948
rect 12980 -4494 13094 -4086
rect 13714 -4494 13876 -4086
rect 15400 -4227 16157 -4186
rect 15400 -4348 15558 -4227
rect 15997 -4348 16157 -4227
rect 15400 -4387 16157 -4348
rect 12980 -4572 13876 -4494
rect 14300 -4744 14624 -4666
rect 14300 -4954 14392 -4744
rect 14550 -4954 14624 -4744
rect 14300 -5036 14624 -4954
rect 10994 -5486 11342 -5446
rect 10994 -5800 11040 -5486
rect 11300 -5800 11342 -5486
rect 10994 -5834 11342 -5800
rect 10216 -6194 10344 -6056
rect -3052 -6518 -2502 -6446
rect -3052 -7126 -2964 -6518
rect -3053 -7204 -2964 -7126
rect -3052 -7226 -2964 -7204
rect -2554 -7126 -2502 -6518
rect 274 -7122 364 -7120
rect 240 -7126 364 -7122
rect -2554 -7156 364 -7126
rect -2554 -7204 286 -7156
rect -2554 -7226 -2502 -7204
rect -3052 -7308 -2502 -7226
rect 274 -7390 286 -7204
rect 354 -7390 364 -7156
rect 274 -7418 364 -7390
rect 2970 -8039 3135 -8005
rect -3048 -8660 -2498 -8572
rect 3101 -8637 3135 -8039
rect -3048 -8696 -2964 -8660
rect -3052 -8788 -2964 -8696
rect -3048 -9368 -2964 -8788
rect -2554 -8696 -2498 -8660
rect 1901 -8671 3135 -8637
rect -2554 -8788 720 -8696
rect -2554 -9368 -2498 -8788
rect 628 -9256 720 -8788
rect 1284 -8978 1664 -8914
rect 1284 -9042 1330 -8978
rect 1618 -9042 1664 -8978
rect 1284 -9066 1664 -9042
rect 1901 -9228 1935 -8671
rect 1812 -9236 1938 -9228
rect 628 -9260 992 -9256
rect 626 -9276 992 -9260
rect 626 -9336 646 -9276
rect 962 -9336 992 -9276
rect 1812 -9290 1832 -9236
rect 1920 -9290 1938 -9236
rect 1812 -9294 1938 -9290
rect 1901 -9295 1935 -9294
rect 626 -9350 992 -9336
rect -3048 -9434 -2498 -9368
rect 420 -9682 1968 -9586
rect 420 -9704 526 -9682
rect -4326 -9892 526 -9704
rect 1804 -9892 1968 -9682
rect -4326 -9940 1968 -9892
rect -4326 -12110 1058 -9940
rect -322 -39220 472 -39194
rect -322 -39290 -276 -39220
rect 422 -39290 472 -39220
rect -322 -39314 472 -39290
rect -1036 -41120 476 -41096
rect -1036 -41188 -260 -41120
rect 424 -41188 476 -41120
rect -1036 -41216 476 -41188
rect -326 -43030 470 -43002
rect -326 -43088 -262 -43030
rect 436 -43088 470 -43030
rect -326 -43118 470 -43088
rect -314 -44940 472 -44906
rect -314 -45004 -284 -44940
rect 436 -45004 472 -44940
rect -314 -45032 472 -45004
rect -324 -46846 488 -46798
rect -324 -46904 -248 -46846
rect 416 -46904 488 -46846
rect -324 -46922 488 -46904
rect -336 -48748 480 -48718
rect -336 -48810 -298 -48748
rect 442 -48810 480 -48748
rect -336 -48836 480 -48810
rect 161022 -80316 166580 -79794
rect 147308 -87889 166580 -80316
rect 132474 -88070 166580 -87889
rect 132474 -88129 148006 -88070
rect 147370 -88143 148000 -88129
rect 10473 -99429 14022 -99129
rect 10473 -100779 10773 -99429
rect 13547 -100779 14022 -99429
rect 10473 -101079 14022 -100779
rect 10583 -105681 14586 -104896
rect 10583 -107252 10989 -105681
rect 13851 -107252 14586 -105681
rect 10583 -107936 14586 -107252
rect -18798 -110928 -12069 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18798 -111995 -12069 -111747
<< via2 >>
rect 62 48122 736 48182
rect 44 46222 766 46280
rect 28 44328 746 44386
rect 78 42418 742 42476
rect 64 40510 738 40566
rect 66 38598 716 38664
rect -2262 33956 -1926 35554
rect -22119 2324 -19207 3207
rect -2468 2398 -1848 3266
rect 3492 2288 4532 3212
rect 811 912 922 1027
rect 8960 5410 10878 6950
rect 8662 2824 8896 3276
rect 12636 3792 13752 4212
rect 148252 3528 151036 3732
rect 15888 3184 16384 3272
rect 10408 1902 10572 2186
rect 14298 2396 14596 2720
rect 15073 2678 15496 2912
rect 7582 260 7642 582
rect 9956 562 10042 698
rect 6880 -556 7024 -472
rect -4990 -1554 -4196 -906
rect 4588 -916 4714 -848
rect 5708 -894 5768 -782
rect 10164 -380 10374 -66
rect 151268 1770 152032 1946
rect 141758 508 143186 868
rect 147540 791 147666 905
rect 150748 68 151082 174
rect 8576 -3338 9764 -2976
rect 7776 -4390 8296 -4148
rect 8224 -4916 9050 -4712
rect 10526 -3898 10794 -3666
rect 14748 -3504 15165 -3198
rect 13094 -4494 13714 -4086
rect 15558 -4348 15997 -4227
rect 14392 -4954 14550 -4744
rect 11040 -5800 11300 -5486
rect 286 -7390 354 -7156
rect 1330 -9042 1618 -8978
rect 526 -9892 1804 -9682
rect -276 -39290 422 -39220
rect -260 -41188 424 -41120
rect -262 -43088 436 -43030
rect -284 -45004 436 -44940
rect -248 -46904 416 -46846
rect -298 -48810 442 -48748
rect 10773 -100779 13547 -99429
rect 10989 -107252 13851 -105681
rect -18327 -111747 -12516 -110928
<< metal3 >>
rect -2 48182 794 48220
rect -2 48122 62 48182
rect 736 48122 794 48182
rect -2 48094 794 48122
rect -2 46280 802 46310
rect -2 46222 44 46280
rect 766 46222 802 46280
rect -2 46192 802 46222
rect 0 44386 800 44412
rect 0 44328 28 44386
rect 746 44328 800 44386
rect 0 44298 800 44328
rect 7474 38032 7928 38152
rect 7808 37496 7928 38032
rect -2200 37376 7928 37496
rect -2200 35752 -2080 37376
rect -2372 35554 -1814 35752
rect -2372 33956 -2262 35554
rect -1926 33956 -1814 35554
rect -2372 33750 -1814 33956
rect -8526 6950 11258 7274
rect -8526 5410 8960 6950
rect 10878 5410 11258 6950
rect -8526 5070 11258 5410
rect -22408 3207 -18497 3481
rect -5176 3446 -2824 3456
rect -5176 3444 -824 3446
rect -22408 2324 -22119 3207
rect -19207 2324 -18497 3207
rect -22408 2088 -18497 2324
rect -5178 3266 -824 3444
rect -5178 3222 -2468 3266
rect -5178 2274 -4942 3222
rect -3104 2398 -2468 3222
rect -1848 2398 -824 3266
rect -3104 2276 -824 2398
rect 3294 3212 4770 3444
rect 3294 2288 3492 3212
rect 4532 2288 4770 3212
rect 8606 3276 8962 3350
rect 8606 2824 8662 3276
rect 8896 2824 8962 3276
rect 8606 2784 8962 2824
rect -3104 2274 706 2276
rect -5178 1392 706 2274
rect 3294 2068 4770 2288
rect 10346 2186 10626 2256
rect 10346 1902 10408 2186
rect 10572 1902 10626 2186
rect 10346 1848 10626 1902
rect -4218 1384 -824 1392
rect -6585 1027 948 1054
rect -6585 912 811 1027
rect 922 912 948 1027
rect -6585 888 948 912
rect 9932 722 10060 730
rect 7552 698 10060 722
rect 7552 582 9956 698
rect 7552 534 7582 582
rect -6584 260 -6152 264
rect -5374 260 1828 264
rect -6584 136 1828 260
rect 7554 260 7582 534
rect 7642 562 9956 582
rect 10042 562 10060 698
rect 7642 536 10060 562
rect 7642 534 9972 536
rect 7642 260 7658 534
rect 7554 234 7658 260
rect 7560 232 7634 234
rect 978 134 1824 136
rect 1636 88 1824 134
rect -6575 30 1086 36
rect -6575 25 1140 30
rect -6575 -98 1191 25
rect -5104 -906 780 -784
rect 1089 -786 1191 -98
rect 1648 -642 1824 88
rect 10076 -66 10462 40
rect 10076 -224 10164 -66
rect 6906 -380 10164 -224
rect 10374 -262 10462 -66
rect 10374 -380 10388 -262
rect 6906 -428 10388 -380
rect 6820 -472 10388 -428
rect 6820 -556 6880 -472
rect 7024 -526 10388 -472
rect 7024 -546 10250 -526
rect 7024 -556 7064 -546
rect 6820 -606 7064 -556
rect 1648 -706 5782 -642
rect 1651 -720 5782 -706
rect 5690 -782 5782 -720
rect 1089 -832 4726 -786
rect 1089 -848 4732 -832
rect 1089 -888 4588 -848
rect -5104 -1554 -4990 -906
rect -4196 -1554 780 -906
rect 4570 -916 4588 -888
rect 4714 -916 4732 -848
rect 5690 -894 5708 -782
rect 5768 -894 5782 -782
rect 5690 -910 5782 -894
rect 4570 -932 4732 -916
rect -5104 -1668 780 -1554
rect -104 -2878 780 -1668
rect 3516 -2650 4164 -2522
rect -104 -3454 916 -2878
rect 8492 -2976 9900 -2888
rect 8492 -3338 8576 -2976
rect 9764 -3338 9900 -2976
rect 8492 -3448 9900 -3338
rect 3728 -3610 4512 -3540
rect 10564 -3600 10851 -3408
rect 3728 -3904 3860 -3610
rect 4402 -3684 4512 -3610
rect 10456 -3666 10854 -3600
rect 10456 -3684 10526 -3666
rect 4402 -3898 10526 -3684
rect 10794 -3898 10854 -3666
rect 4402 -3904 10854 -3898
rect 3728 -3966 10854 -3904
rect 3728 -3972 10852 -3966
rect 7680 -4148 8400 -4072
rect 7680 -4390 7776 -4148
rect 8296 -4390 8400 -4148
rect 7680 -4456 8400 -4390
rect 8118 -4712 9202 -4628
rect 8118 -4916 8224 -4712
rect 9050 -4916 9202 -4712
rect 8118 -4990 9202 -4916
rect 274 -7122 364 -7120
rect 240 -7156 364 -7122
rect 240 -7202 286 -7156
rect 274 -7390 286 -7202
rect 354 -7390 364 -7156
rect 274 -7418 364 -7390
rect 274 -8822 342 -7418
rect 274 -8890 3124 -8822
rect 1284 -8978 1666 -8954
rect 1284 -9042 1330 -8978
rect 1618 -9042 1666 -8978
rect 1284 -9066 1666 -9042
rect 8206 -9146 9262 -9048
rect 8206 -9532 8304 -9146
rect 9182 -9532 9262 -9146
rect 420 -9682 1968 -9586
rect 8206 -9596 9262 -9532
rect 420 -9892 526 -9682
rect 1804 -9892 1968 -9682
rect 420 -9940 1968 -9892
rect 10564 -10166 10851 -3972
rect 10994 -5486 11342 -5446
rect 10994 -5800 11040 -5486
rect 11300 -5800 11342 -5486
rect 10994 -5834 11342 -5800
rect -11764 -11810 10786 -10166
rect 9785 -30482 11338 -30481
rect 11530 -30482 12425 30261
rect 12520 4212 13874 4286
rect 12520 3792 12636 4212
rect 13752 3792 13874 4212
rect 12520 3712 13874 3792
rect 15833 3272 16452 3314
rect 15833 3184 15888 3272
rect 16384 3184 16452 3272
rect 15833 3149 16452 3184
rect 14983 2912 15595 2991
rect 14236 2735 14374 2792
rect 14482 2735 14682 2792
rect 14236 2720 14682 2735
rect 14236 2396 14298 2720
rect 14596 2396 14682 2720
rect 14983 2678 15073 2912
rect 15496 2678 15595 2912
rect 14983 2604 15595 2678
rect 14236 2318 14682 2396
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 141714 440 143268 508
rect 147523 905 147705 6789
rect 148146 3732 151160 3818
rect 148146 3528 148252 3732
rect 151036 3528 151160 3732
rect 148146 3436 151160 3528
rect 151204 1946 152196 2020
rect 151204 1770 151268 1946
rect 152032 1770 152196 1946
rect 151204 1725 152196 1770
rect 147523 791 147540 905
rect 147666 791 147705 905
rect 142650 232 143030 440
rect 147523 232 147705 791
rect 142650 174 151159 232
rect 142650 68 150748 174
rect 151082 68 151159 174
rect 142650 50 151159 68
rect 142650 -140 143030 50
rect 15062 -520 147620 -140
rect 142551 -1206 144558 -1108
rect 151336 -1204 151438 -1014
rect 149920 -1206 151438 -1204
rect 142264 -1210 151438 -1206
rect 142264 -1410 142634 -1210
rect 144396 -1310 151438 -1210
rect 144396 -1410 151378 -1310
rect 142264 -1502 151378 -1410
rect 14666 -3198 15268 -3130
rect 14666 -3504 14748 -3198
rect 15165 -3504 15268 -3198
rect 14666 -3599 15268 -3504
rect 12980 -4086 13876 -3948
rect 12980 -4494 13094 -4086
rect 13714 -4494 13876 -4086
rect 15400 -4227 16157 -4186
rect 15400 -4348 15558 -4227
rect 15997 -4348 16157 -4227
rect 15400 -4387 16157 -4348
rect 12980 -4572 13876 -4494
rect 14300 -4744 14624 -4666
rect 14300 -4954 14392 -4744
rect 14550 -4954 14624 -4744
rect 14300 -5036 14624 -4954
rect 9785 -31539 12425 -30482
rect 9785 -33235 10843 -31539
rect -322 -39220 472 -39194
rect -322 -39290 -276 -39220
rect 422 -39290 472 -39220
rect -322 -39314 472 -39290
rect -320 -41120 482 -41092
rect -320 -41188 -260 -41120
rect 424 -41188 482 -41120
rect -320 -41212 482 -41188
rect -12084 -95510 10770 -87288
rect 10473 -99429 14022 -99129
rect 10473 -100779 10773 -99429
rect 13547 -100779 14022 -99429
rect 10473 -101079 14022 -100779
rect 10583 -105681 14586 -104896
rect 10583 -107252 10989 -105681
rect 13851 -107252 14586 -105681
rect 10583 -107936 14586 -107252
rect -18798 -110928 -12069 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18798 -111995 -12069 -111747
<< via3 >>
rect -22119 2324 -19207 3207
rect -4942 2274 -3104 3222
rect -2468 2398 -1848 3266
rect 3492 2288 4532 3212
rect 8662 2824 8896 3276
rect 10408 1902 10572 2186
rect -4990 -1554 -4196 -906
rect 8576 -3338 9764 -2976
rect 3860 -3904 4402 -3610
rect 7776 -4390 8296 -4148
rect 8224 -4916 9050 -4712
rect 1330 -9042 1618 -8978
rect 8304 -9532 9182 -9146
rect 526 -9892 1804 -9682
rect 11040 -5800 11300 -5486
rect 12636 3792 13752 4212
rect 14298 2396 14596 2720
rect 15073 2678 15496 2912
rect 141758 508 143186 868
rect 148252 3528 151036 3732
rect 151268 1770 152032 1946
rect 142634 -1410 144396 -1210
rect 14748 -3504 15165 -3198
rect 13094 -4494 13714 -4086
rect 15558 -4348 15997 -4227
rect 14392 -4954 14550 -4744
rect 10773 -100779 13547 -99429
rect 10989 -107252 13851 -105681
rect -18327 -111747 -12516 -110928
<< metal4 >>
rect -42087 103024 17476 108254
rect -42087 98072 17648 103024
rect 16921 94385 17619 98072
rect -4264 4744 890 7690
rect -22408 3207 -18497 3481
rect -22408 2324 -22119 3207
rect -19207 2324 -18497 3207
rect -22408 2088 -18497 2324
rect -5176 3222 -2824 3456
rect -5176 2274 -4942 3222
rect -3104 2274 -2824 3222
rect -5176 2076 -2824 2274
rect -2626 3266 -1628 4744
rect 12492 4212 13874 4296
rect 12492 3792 12636 4212
rect 13752 3792 13874 4212
rect 12492 3714 13874 3792
rect -2626 2398 -2468 3266
rect -1848 2398 -1628 3266
rect -2626 2132 -1628 2398
rect 3294 3212 4770 3444
rect 3294 2288 3492 3212
rect 4532 2288 4770 3212
rect 8606 3278 8962 3350
rect 8606 2824 8654 3278
rect 8910 2824 8962 3278
rect 8606 2784 8962 2824
rect 14983 2922 15595 2991
rect 14276 2788 14374 2794
rect 3294 2068 4770 2288
rect 14238 2735 14374 2788
rect 14482 2735 14683 2794
rect 14238 2720 14683 2735
rect 14238 2396 14298 2720
rect 14596 2692 14683 2720
rect 14596 2396 14684 2692
rect 14983 2674 15073 2922
rect 15499 2674 15595 2922
rect 14983 2604 15595 2674
rect 14238 2252 14684 2396
rect 9102 2186 14684 2252
rect 9102 1902 10408 2186
rect 10572 1902 14684 2186
rect 9102 1844 14684 1902
rect -5190 -682 1060 1212
rect 10930 128 11338 1844
rect 13472 1692 14040 1844
rect 15722 1692 16290 4472
rect 13472 1124 14206 1692
rect 14808 1124 16290 1692
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 141714 440 143268 508
rect 140356 128 141376 178
rect -5108 -906 -4096 -682
rect -5108 -1554 -4990 -906
rect -4196 -1554 -4096 -906
rect -5108 -1672 -4096 -1554
rect 10930 -866 141618 128
rect -10346 -4062 -4938 -3018
rect 3728 -3540 4490 -2808
rect 8492 -2976 9900 -2888
rect 8492 -3338 8576 -2976
rect 9764 -3338 9900 -2976
rect 8492 -3448 9900 -3338
rect 3728 -3610 4512 -3540
rect 3728 -3904 3860 -3610
rect 4402 -3904 4512 -3610
rect 3728 -3972 4512 -3904
rect 5716 -4062 6490 -4032
rect 10930 -4062 11338 -866
rect 140268 -870 141376 -866
rect 140268 -1102 141272 -870
rect 140268 -1210 144598 -1102
rect 140268 -1410 142634 -1210
rect 144396 -1410 144598 -1210
rect 140268 -1492 144598 -1410
rect 14666 -3198 15268 -3130
rect 14666 -3504 14748 -3198
rect 15165 -3504 15268 -3198
rect 14666 -3599 15268 -3504
rect -10346 -4148 11338 -4062
rect -10346 -4390 7776 -4148
rect 8296 -4390 11338 -4148
rect -10346 -4470 11338 -4390
rect -10346 -4950 -4938 -4470
rect 324 -8660 732 -4470
rect 5026 -4472 5434 -4470
rect 5026 -5688 5434 -5608
rect 5716 -5828 6490 -4470
rect 8118 -4712 9202 -4628
rect 8118 -4916 8224 -4712
rect 9050 -4766 9202 -4712
rect 10930 -4630 11338 -4470
rect 12980 -4086 13876 -3948
rect 12980 -4494 13094 -4086
rect 13714 -4494 13876 -4086
rect 15400 -4227 16157 -4186
rect 15400 -4348 15558 -4227
rect 15997 -4348 16157 -4227
rect 15400 -4387 16157 -4348
rect 12980 -4572 13876 -4494
rect 10930 -4666 11342 -4630
rect 10930 -4744 14628 -4666
rect 9050 -4866 9544 -4766
rect 9050 -4916 9202 -4866
rect 8118 -4990 9202 -4916
rect 9444 -7094 9544 -4866
rect 10930 -4954 14392 -4744
rect 14550 -4954 14628 -4744
rect 10930 -5038 14628 -4954
rect 10930 -5432 11338 -5038
rect 10378 -5486 11338 -5432
rect 10378 -5800 11040 -5486
rect 11300 -5800 11338 -5486
rect 10378 -5840 11338 -5800
rect 145536 -7134 146104 4496
rect 148146 3732 151152 4574
rect 148146 3528 148252 3732
rect 151036 3528 151152 3732
rect 148146 3436 151152 3528
rect 151204 1946 152196 2020
rect 151204 1770 151268 1946
rect 152032 1770 152196 1946
rect 151204 1725 152196 1770
rect 151204 -700 151550 1725
rect 324 -8978 1666 -8660
rect 324 -9042 1330 -8978
rect 1618 -9042 1666 -8978
rect 324 -9068 1666 -9042
rect 8206 -9146 9432 -9052
rect 8206 -9532 8304 -9146
rect 9182 -9532 9432 -9146
rect 420 -9682 1968 -9586
rect 8206 -9592 9432 -9532
rect 420 -9704 526 -9682
rect -4326 -9892 526 -9704
rect 1804 -9892 1968 -9682
rect -4326 -9940 1968 -9892
rect -4326 -12110 1058 -9940
rect 10473 -99429 14022 -99129
rect 10473 -100779 10773 -99429
rect 13547 -100779 14022 -99429
rect 10473 -101079 14022 -100779
rect 10583 -105681 14586 -104896
rect 10583 -107252 10989 -105681
rect 13851 -107252 14586 -105681
rect 10583 -107936 14586 -107252
rect -18798 -110928 -12069 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18798 -111995 -12069 -111747
rect -12432 -113425 -6589 -112623
rect -12432 -114424 -11561 -113425
rect -13282 -114761 -11561 -114424
rect -12432 -115281 -11561 -114761
rect -7941 -115281 -6589 -113425
rect -12432 -116014 -6589 -115281
<< via4 >>
rect -22119 2324 -19207 3207
rect -4942 2274 -3104 3222
rect 12636 3792 13752 4212
rect -2468 2398 -1848 3266
rect 3492 2288 4532 3212
rect 8654 3276 8910 3278
rect 8654 2824 8662 3276
rect 8662 2824 8896 3276
rect 8896 2824 8910 3276
rect 15073 2912 15499 2922
rect 15073 2678 15496 2912
rect 15496 2678 15499 2912
rect 15073 2674 15499 2678
rect 141758 508 143186 868
rect 8576 -3338 9764 -2976
rect 14748 -3504 15165 -3198
rect 13094 -4494 13714 -4086
rect 8322 -9526 9176 -9146
rect 10773 -100779 13547 -99429
rect 10989 -107252 13851 -105681
rect -18327 -111747 -12516 -110928
rect -11561 -115281 -7941 -113425
<< metal5 >>
rect 146169 5724 146682 5849
rect 12502 4212 13877 4293
rect 12502 3792 12636 4212
rect 13752 3792 13877 4212
rect -22408 3463 -18497 3481
rect 12502 3463 13877 3792
rect -22408 3278 13877 3463
rect -22408 3266 8654 3278
rect -22408 3222 -2468 3266
rect -22408 3207 -4942 3222
rect -22408 2324 -22119 3207
rect -19207 2324 -4942 3207
rect -22408 2274 -4942 2324
rect -3104 2398 -2468 3222
rect -1848 3212 8654 3266
rect -1848 2398 3492 3212
rect -3104 2288 3492 2398
rect 4532 2824 8654 3212
rect 8910 2824 13877 3278
rect 4532 2288 13877 2824
rect 14983 2922 15595 2991
rect 14983 2674 15073 2922
rect 15499 2674 15595 2922
rect 14983 2604 15595 2674
rect -3104 2274 13877 2288
rect 15585 2276 15595 2604
rect -22408 2088 13877 2274
rect 3294 2068 4770 2088
rect 8483 -2702 9858 2088
rect 141714 944 143268 950
rect 138862 868 143292 944
rect 138862 508 141758 868
rect 143186 508 143292 868
rect 138862 442 143292 508
rect 13033 82 13831 297
rect 138874 82 140192 442
rect 141714 440 143268 442
rect 13033 -786 141618 82
rect 8480 -2726 9860 -2702
rect 13033 -2726 13831 -786
rect 138874 -852 140192 -786
rect 8458 -2976 13866 -2726
rect 8458 -3338 8576 -2976
rect 9764 -3338 13866 -2976
rect 8458 -3524 13866 -3338
rect 8480 -3640 9860 -3524
rect 10411 -8791 11209 -3524
rect 12983 -4086 13866 -3524
rect 12983 -4494 13094 -4086
rect 13714 -4494 13866 -4086
rect 12983 -4559 13866 -4494
rect 12983 -4565 13781 -4559
rect 146169 -7895 146759 5724
rect 8987 -9052 11209 -8791
rect 8206 -9146 11209 -9052
rect 8206 -9526 8322 -9146
rect 9176 -9526 11209 -9146
rect 8206 -9589 11209 -9526
rect 8206 -9592 9432 -9589
rect 15603 -98230 16321 -97802
rect -12568 -99429 16452 -98230
rect -12568 -100779 10773 -99429
rect 13547 -100779 16452 -99429
rect -12568 -105681 16452 -100779
rect -12568 -107252 10989 -105681
rect 13851 -107252 16452 -105681
rect -12568 -109101 16452 -107252
rect -12596 -110641 16511 -109101
rect -18778 -110654 16511 -110641
rect -18798 -110928 16511 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 16511 -110928
rect -18798 -111995 16511 -111747
rect -18778 -112016 16511 -111995
rect -12596 -113425 16511 -112016
rect -12596 -115281 -11561 -113425
rect -7941 -115281 16511 -113425
rect -12596 -116321 16511 -115281
use cmfb_pmos  cmfb_pmos_0
timestamp 1727004346
transform 1 0 148450 0 1 -716
box -158 762 4965 2374
use comparator_final_compact  comparator_final_compact_0
timestamp 1727642364
transform -1 0 9078 0 1 -7110
box -2532 -2214 8345 1614
use full_stage_modified  full_stage_modified_0
timestamp 1727007906
transform 1 0 3520 0 1 -3410
box 8 8 4397 4640
use reconfigurable_CP  reconfigurable_CP_0
timestamp 1727647182
transform 1 0 16242 0 -1 63194
box -16242 -34774 130792 69994
use reconfigurable_CP  reconfigurable_CP_1
timestamp 1727647182
transform 1 0 15920 0 1 -63814
box -16242 -34774 130792 69994
use reference0_9  reference0_9_0
timestamp 1699232519
transform 0 -1 151950 1 0 -1600
box -66 -1120 1022 620
use reference  reference_1
timestamp 1727087973
transform 0 1 9868 -1 0 4356
box -32 -858 1828 500
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_0
timestamp 1699146224
transform -1 0 150592 0 -1 7074
box -3186 -3040 3186 3040
use sky130_fd_pr__nfet_01v8_PXJ6TW  sky130_fd_pr__nfet_01v8_PXJ6TW_0
timestamp 1699271609
transform 1 0 148196 0 1 1206
box -108 -126 108 126
use sky130_fd_pr__nfet_01v8_PXJ6TW  sky130_fd_pr__nfet_01v8_PXJ6TW_1
timestamp 1699271609
transform 1 0 148198 0 1 446
box -108 -126 108 126
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1693170804
transform -1 0 1322 0 1 -9508
box -38 -48 314 592
use source_follower_buffer  source_follower_buffer_0
timestamp 1726987743
transform 1 0 14893 0 1 -4323
box -657 184 577 768
use source_follower_buffer  source_follower_buffer_1
timestamp 1726987743
transform 1 0 14975 0 -1 3723
box -657 184 577 768
<< labels >>
flabel metal5 15603 -105367 15617 -105363 0 FreeSans 4800 90 0 0 digital_gnd
flabel metal4 16921 102321 17619 103019 0 FreeSans 4800 90 0 0 digital_vdd
flabel space 8228 39660 9060 39802 0 FreeSans 3200 0 0 0 scan_out
flabel space 148376 1942 148438 2082 0 FreeSans 2400 90 0 0 vd1
flabel space 148306 -658 148460 -292 0 FreeSans 2400 90 0 0 vd2
flabel metal4 -30725 98072 -20543 108254 0 FreeSans 16000 0 0 0 digital_vdd_1.8V
flabel space -6158 -95630 2366 -87288 0 FreeSans 16000 0 0 0 clock(internal)_50MHz
flabel metal5 -6522 -108146 -1140 -101858 0 FreeSans 16000 0 0 0 Digital_gnd
flabel metal2 157929 79019 166338 87428 0 FreeSans 16000 0 0 0 vout+
flabel metal2 153340 2296 153890 2902 0 FreeSans 8000 0 0 0 vd1
flabel space 153456 -2960 154006 -2354 0 FreeSans 8000 0 0 0 vd2
flabel space 153424 -88070 161700 -79794 0 FreeSans 16000 0 0 0 vout-
flabel space -6574 46716 -5648 48142 0 FreeSans 8000 0 0 0 clk_external
flabel metal2 -7251 42824 -5689 44386 0 FreeSans 8000 0 0 0 scan_in
flabel metal2 -8468 40388 -6658 42012 0 FreeSans 8000 0 0 0 scan_en
flabel metal2 -8260 38108 -6042 39556 0 FreeSans 8000 0 0 0 reset
flabel space -5816 -100 -5606 34 0 FreeSans 1600 0 0 0 drain1
flabel space -5822 136 -5612 270 0 FreeSans 1600 0 0 0 drain2
flabel space -5812 1068 -5638 1152 0 FreeSans 1600 0 0 0 ib2_1uA
flabel psubdiff -11610 -11898 -9966 -10254 0 FreeSans 8000 0 0 0 v_int-
flabel metal3 -8526 5070 -6322 7274 0 FreeSans 8000 0 0 0 v_int+
flabel space -10456 2110 -8262 3522 0 FreeSans 6400 0 0 0 analog_gnd
flabel metal4 -10346 -4950 -8000 -3018 0 FreeSans 6400 0 0 0 analog_vdd_1.8V
rlabel via1 912 962 912 962 1 ib2
flabel space 6446 -38882 7520 -38354 0 FreeSans 4800 0 0 0 scan_out
<< end >>
