* SPICE3 file created from reconfigurable_CP1.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_HRDN5X a_n129_n130# a_n369_n42# a_543_64# a_63_n130#
+ a_159_64# a_n417_64# a_687_n42# a_303_n42# a_n561_n42# a_n321_n130# a_n749_n42#
+ a_639_n130# a_n81_n42# a_399_n42# a_n273_n42# a_15_n42# a_447_n130# a_n609_64# a_591_n42#
+ a_207_n42# a_n465_n42# a_351_64# a_255_n130# a_n33_64# a_n225_64# a_n705_n130# a_n177_n42#
+ a_n657_n42# a_495_n42# a_111_n42# a_n513_n130# VSUBS
X0 a_303_n42# a_255_n130# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_591_n42# a_543_64# a_495_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_207_n42# a_159_64# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_399_n42# a_351_64# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_495_n42# a_447_n130# a_399_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_687_n42# a_639_n130# a_591_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n561_n42# a_n609_64# a_n657_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n657_n42# a_n705_n130# a_n749_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X8 a_n465_n42# a_n513_n130# a_n561_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n369_n42# a_n417_64# a_n465_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n273_n42# a_n321_n130# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n81_n42# a_n129_n130# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n177_n42# a_n225_64# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MH6KF8 c1_n1046_n900# m3_n1086_n940# VSUBS
X0 c1_n1046_n900# m3_n1086_n940# sky130_fd_pr__cap_mim_m3_1 l=9 w=9
C0 m3_n1086_n940# c1_n1046_n900# 7.77654f
C1 m3_n1086_n940# VSUBS 3.30833f
.ends

.subckt nmos_dnw3 vin out1 out2 clk clkb vs VSUBS
X0 clkb clk vin vs sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.126 ps=1.44 w=0.42 l=0.15
X1 vin clkb clk vs sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.1302 ps=1.46 w=0.42 l=0.15
X2 out2 clk vin vs sky130_fd_pr__nfet_01v8 ad=1.65 pd=7.1 as=0.945 ps=3.63 w=3 l=1
X3 vin clkb out1 vs sky130_fd_pr__nfet_01v8 ad=0.945 pd=3.63 as=1.65 ps=7.1 w=3 l=1
C0 vs VSUBS 6.63893f
.ends

.subckt sky130_fd_pr__pfet_01v8_FBZ64Q a_n81_n126# a_399_n126# a_351_n223# a_n417_n223#
+ a_207_n126# a_n225_n223# a_n461_n126# a_n369_n126# a_63_157# a_303_n126# a_255_157#
+ a_n33_n223# a_15_n126# a_n177_n126# a_n129_157# a_111_n126# w_n497_n226# a_n273_n126#
+ a_159_n223# a_n321_157# VSUBS
X0 a_n273_n126# a_n321_157# a_n369_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 a_207_n126# a_159_n223# a_111_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X2 a_n177_n126# a_n225_n223# a_n273_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 a_111_n126# a_63_157# a_15_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_399_n126# a_351_n223# a_303_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_n81_n126# a_n129_157# a_n177_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X6 a_15_n126# a_n33_n223# a_n81_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X7 a_n369_n126# a_n417_n223# a_n461_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X8 a_303_n126# a_255_157# a_207_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_5ACVEW a_n129_n130# a_63_n130# a_n81_n42# a_15_n42#
+ a_n173_n42# a_n33_64# a_111_n42# VSUBS
X0 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n81_n42# a_n129_n130# a_n173_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGLN5 a_n129_n130# a_n369_n42# a_1215_n130# a_543_64#
+ a_63_n130# a_159_64# a_n1089_n130# a_n849_n42# a_n417_64# a_n801_64# a_687_n42#
+ a_303_n42# a_1167_n42# a_n561_n42# a_n321_n130# a_n1041_n42# a_639_n130# a_n1185_64#
+ a_1023_n130# a_n1281_n130# a_n81_n42# a_399_n42# a_879_n42# a_n273_n42# a_735_64#
+ a_n753_n42# a_15_n42# a_n897_n130# a_n1233_n42# a_831_n130# a_447_n130# a_n609_64#
+ a_1071_n42# a_591_n42# a_1119_64# a_n993_64# a_207_n42# a_n465_n42# a_n945_n42#
+ a_351_64# a_783_n42# a_255_n130# a_n33_64# a_n225_64# a_n705_n130# a_1263_n42# a_927_64#
+ a_n177_n42# a_n657_n42# a_n1325_n42# a_n1137_n42# a_495_n42# a_111_n42# a_975_n42#
+ a_n513_n130# VSUBS
X0 a_303_n42# a_255_n130# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_591_n42# a_543_64# a_495_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_207_n42# a_159_64# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_399_n42# a_351_64# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_495_n42# a_447_n130# a_399_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_687_n42# a_639_n130# a_591_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_783_n42# a_735_64# a_687_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_975_n42# a_927_64# a_879_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n1041_n42# a_n1089_n130# a_n1137_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_879_n42# a_831_n130# a_783_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n1233_n42# a_n1281_n130# a_n1325_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X11 a_n1137_n42# a_n1185_64# a_n1233_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n561_n42# a_n609_64# a_n657_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1071_n42# a_1023_n130# a_975_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1263_n42# a_1215_n130# a_1167_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n945_n42# a_n993_64# a_n1041_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n753_n42# a_n801_64# a_n849_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n657_n42# a_n705_n130# a_n753_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n465_n42# a_n513_n130# a_n561_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n369_n42# a_n417_64# a_n465_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_1167_n42# a_1119_64# a_1071_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n849_n42# a_n897_n130# a_n945_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n273_n42# a_n321_n130# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n81_n42# a_n129_n130# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n177_n42# a_n225_64# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_VR4B8J a_1119_157# a_783_n126# a_n81_n126# a_n849_n126#
+ a_399_n126# a_n1041_n126# a_351_157# a_495_n126# a_n945_n126# a_n33_157# a_n129_n223#
+ a_n513_n223# a_1215_n223# a_63_n223# a_n1089_n223# a_n225_157# a_591_n126# a_n657_n126#
+ a_207_n126# a_543_157# a_n1325_n126# a_n369_n126# a_n753_n126# a_n321_n223# a_303_n126#
+ a_1023_n223# a_639_n223# a_n1281_n223# a_n417_157# a_n465_n126# a_1167_n126# a_735_157#
+ a_15_n126# a_n561_n126# a_n993_157# a_n177_n126# a_n897_n223# w_n1361_n226# a_1263_n126#
+ a_879_n126# a_111_n126# a_831_n223# a_n609_157# a_447_n223# a_n273_n126# a_n1137_n126#
+ a_975_n126# a_927_157# a_n1185_157# a_n1233_n126# a_n801_157# a_1071_n126# a_687_n126#
+ a_255_n223# a_n705_n223# a_159_157# VSUBS
X0 a_n273_n126# a_n321_n223# a_n369_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 a_n1233_n126# a_n1281_n223# a_n1325_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X2 a_591_n126# a_543_157# a_495_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 a_n849_n126# a_n897_n223# a_n945_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_207_n126# a_159_157# a_111_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_n177_n126# a_n225_157# a_n273_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X6 a_n1137_n126# a_n1185_157# a_n1233_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X7 a_495_n126# a_447_n223# a_399_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X8 a_n561_n126# a_n609_157# a_n657_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X9 a_111_n126# a_63_n223# a_15_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X10 a_783_n126# a_735_157# a_687_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X11 a_1071_n126# a_1023_n223# a_975_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X12 a_399_n126# a_351_157# a_303_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X13 a_n465_n126# a_n513_n223# a_n561_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X14 a_687_n126# a_639_n223# a_591_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X15 a_n753_n126# a_n801_157# a_n849_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X16 a_975_n126# a_927_157# a_879_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X17 a_n81_n126# a_n129_n223# a_n177_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X18 a_15_n126# a_n33_157# a_n81_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X19 a_1263_n126# a_1215_n223# a_1167_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X20 a_n1041_n126# a_n1089_n223# a_n1137_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X21 a_n369_n126# a_n417_157# a_n465_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X22 a_n657_n126# a_n705_n223# a_n753_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X23 a_879_n126# a_831_n223# a_783_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X24 a_n945_n126# a_n993_157# a_n1041_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X25 a_1167_n126# a_1119_157# a_1071_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X26 a_303_n126# a_255_n223# a_207_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
C0 w_n1361_n226# VSUBS 3.66914f
.ends

.subckt inverter_27x m1_n804_1398# m1_540_1398# m1_156_1398# m1_n36_1398# m1_732_1398#
+ m1_n1102_1398# m1_348_1398# m1_n1188_1398# m1_n996_1398# m1_n228_1398# m1_n1188_1912#
+ m1_924_1398# m1_1309_1398# a_n1158_1658# m1_n420_1398# m1_1116_1398# w_1358_2036#
+ m1_n612_1398# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1658# m1_n228_1398# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# a_n1158_1658# a_n1158_1658#
+ m1_n1102_1398# m1_n1102_1398# m1_1309_1398# m1_n420_1398# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_540_1398#
+ m1_n1102_1398# m1_n1102_1398# a_n1158_1658# m1_n612_1398# m1_156_1398# a_n1158_1658#
+ m1_n1102_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_732_1398#
+ a_n1158_1658# a_n1158_1658# m1_348_1398# m1_n1102_1398# m1_n804_1398# a_n1158_1658#
+ m1_924_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# m1_n36_1398# m1_n1102_1398# m1_n1188_1398# m1_n996_1398# m1_n1102_1398#
+ m1_n1102_1398# m1_1116_1398# a_n1158_1658# VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1658# m1_n1188_1912# m1_1309_1398# m1_1309_1398#
+ m1_n1188_1912# m1_1309_1398# a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ m1_n1188_1912# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ a_n1158_1658# m1_n1188_1912# a_n1158_1658# w_1358_2036# m1_1309_1398# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_1309_1398# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# a_n1158_1658# m1_1309_1398# a_n1158_1658# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
C0 a_n1158_1658# VSUBS 6.394793f
C1 w_1358_2036# VSUBS 3.688076f
.ends

.subckt sky130_fd_pr__nfet_01v8_KMMFCM a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_29EZRJ a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_FL984Q a_n81_n126# a_n33_157# a_n129_n223# a_63_n223#
+ a_n173_n126# a_15_n126# a_111_n126# w_n209_n226# VSUBS
X0 a_111_n126# a_63_n223# a_15_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 a_n81_n126# a_n129_n223# a_n173_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X2 a_15_n126# a_n33_157# a_n81_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_FXZ64Q a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_D4CDWR a_n369_n42# a_n225_n130# a_303_n42# a_n81_n42#
+ a_399_n42# a_n33_n130# a_n273_n42# a_n461_n42# a_15_n42# a_n321_64# a_207_n42# a_159_n130#
+ a_n177_n42# a_351_n130# a_255_64# a_n417_n130# a_111_n42# a_n129_64# a_63_64# VSUBS
X0 a_303_n42# a_255_64# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_207_n42# a_159_n130# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_399_n42# a_351_n130# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n369_n42# a_n417_n130# a_n461_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4 a_15_n42# a_n33_n130# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_111_n42# a_63_64# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n273_n42# a_n321_64# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n81_n42# a_n129_64# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n177_n42# a_n225_n130# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_DQBD8A a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt clock clk_in vdd gnd clk clkb
Xsky130_fd_pr__pfet_01v8_FBZ64Q_0 vdd a_3246_118# a_2402_572# a_2402_572# a_3246_118#
+ a_2402_572# vdd a_3246_118# a_2402_572# vdd a_2402_572# a_2402_572# a_3246_118#
+ a_3246_118# a_2402_572# vdd vdd vdd a_2402_572# a_2402_572# gnd sky130_fd_pr__pfet_01v8_FBZ64Q
Xsky130_fd_pr__nfet_01v8_5ACVEW_0 a_344_n986# a_344_n986# a_2402_572# gnd gnd a_344_n986#
+ a_2402_572# gnd sky130_fd_pr__nfet_01v8_5ACVEW
Xinverter_27x_0 clk clk clk clk clk gnd clk clk clk clk vdd clk clk a_3246_118# clk
+ clk vdd clk gnd inverter_27x
Xsky130_fd_pr__nfet_01v8_KMMFCM_0 a_134_122# clk_in gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_1 a_416_120# a_344_102# sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42#
+ gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_2 sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42# a_134_122#
+ gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__pfet_01v8_29EZRJ_0 vdd vdd a_134_122# clk_in gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FL984Q_0 a_2402_572# a_344_n986# a_344_n986# a_344_n986#
+ vdd vdd a_2402_572# vdd gnd sky130_fd_pr__pfet_01v8_FL984Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 vdd vdd a_1230_122# m1_998_498# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_1 a_416_120# vdd vdd a_344_102# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 vdd vdd a_1430_122# a_1230_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_2 vdd vdd a_416_120# a_134_122# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_2 vdd vdd a_344_n986# a_1430_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_3 vdd vdd m1_998_498# a_786_n2# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__nfet_01v8_D4CDWR_0 a_3246_118# a_2402_572# gnd gnd a_3246_118# a_2402_572#
+ gnd gnd a_3246_118# a_2402_572# a_3246_118# a_2402_572# a_3246_118# a_2402_572#
+ a_2402_572# a_2402_572# gnd a_2402_572# a_2402_572# gnd sky130_fd_pr__nfet_01v8_D4CDWR
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 m1_998_498# a_786_n2# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 a_1230_122# m1_998_498# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_2 a_1430_122# a_1230_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_3 a_344_n986# a_1430_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
X0 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X2 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 vdd a_344_102# a_2020_n482# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X7 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X9 a_786_n912# a_586_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X10 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X11 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X12 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X13 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X17 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X20 a_286_n478# clk_in gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.15
X21 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X22 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X24 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_586_n2# a_416_120# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X27 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X28 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X30 a_786_n912# a_586_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X31 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X32 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 vdd a_344_n986# a_286_n960# vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.1827 ps=1.55 w=1.26 l=0.15
X34 a_344_102# a_1394_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X35 a_992_n918# a_786_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X36 a_1192_n918# a_992_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X37 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X38 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X39 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1394_n918# a_1192_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X42 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X43 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X46 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X48 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X49 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X51 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X52 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_586_n912# a_286_n960# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X54 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X55 a_586_n2# a_416_120# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X56 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X57 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X58 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X59 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X61 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X63 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X66 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X68 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_786_n2# a_586_n2# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X72 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_286_n960# clk_in vdd vdd sky130_fd_pr__pfet_01v8 ad=0.1827 pd=1.55 as=0.3654 ps=3.1 w=1.26 l=0.15
X74 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X75 a_286_n960# a_344_n986# a_286_n478# gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.15
X76 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X77 a_586_n912# a_286_n960# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X78 a_1394_n918# a_1192_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X79 a_1192_n918# a_992_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X80 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X81 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X82 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X83 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X84 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X85 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X86 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X87 a_344_102# a_1394_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X88 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X89 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X90 gnd a_344_102# a_2020_n482# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X91 a_992_n918# a_786_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X92 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X93 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X94 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X95 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X96 a_786_n2# a_586_n2# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X97 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
C0 a_2432_n962# vdd 7.043292f
C1 a_2432_n962# clkb 2.67187f
C2 a_2020_n482# vdd 2.656852f
C3 clkb vdd 7.306418f
C4 clkb gnd 5.097592f
C5 a_2432_n962# gnd 8.705547f
C6 a_2020_n482# gnd 2.565399f
C7 vdd gnd 26.103016f
C8 a_344_102# gnd 2.811321f
C9 a_2402_572# gnd 2.314155f
C10 a_344_n986# gnd 2.426004f
C11 a_3246_118# gnd 6.789812f
.ends

.subckt buffer_digital i in VDD GND
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 VDD VDD a_116_148# i GND sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 VDD VDD in a_116_148# GND sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 a_116_148# i GND GND sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 in a_116_148# GND GND sky130_fd_pr__nfet_01v8_DQBD8A
.ends

.subckt sky130_fd_pr__pfet_01v8_4ZKXAA a_63_n42# a_n417_n42# a_303_n139# w_n545_n142#
+ a_255_n42# a_n465_n139# a_n129_n42# a_111_n139# a_447_n42# a_n273_n139# a_n177_73#
+ a_n321_n42# a_207_73# a_n509_n42# a_159_n42# a_15_73# a_n81_n139# a_351_n42# a_n33_n42#
+ a_n369_73# a_n225_n42# a_399_73# VSUBS
X0 a_n33_n42# a_n81_n139# a_n129_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_351_n42# a_303_n139# a_255_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n139# a_63_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_73# a_159_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_447_n42# a_399_73# a_351_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_73# a_n417_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n225_n42# a_n273_n139# a_n321_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n139# a_n509_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X8 a_n129_n42# a_n177_73# a_n225_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_63_n42# a_15_73# a_n33_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_9LGCGE a_15_n130# a_n561_n130# a_63_n42# a_n989_n42#
+ a_n177_n130# a_n417_n42# a_n465_64# a_255_n42# a_495_64# a_735_n42# a_n129_n42#
+ a_n609_n42# a_111_64# a_447_n42# a_927_n42# a_783_n130# a_n321_n42# a_399_n130#
+ a_n657_64# a_n801_n42# a_687_64# a_n945_n130# a_159_n42# a_639_n42# a_n513_n42#
+ a_n897_n42# a_591_n130# a_n81_64# a_n273_64# a_351_n42# a_207_n130# a_303_64# a_n33_n42#
+ a_831_n42# a_n369_n130# a_n753_n130# a_n849_64# a_n225_n42# a_n705_n42# a_879_64#
+ a_543_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n897_n42# a_n945_n130# a_n989_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_49FP49 a_63_n42# a_n989_n42# a_n369_n139# a_n753_n139#
+ a_n417_n42# a_687_73# w_n1025_n142# a_255_n42# a_735_n42# a_n81_73# a_n273_73# a_n129_n42#
+ a_15_n139# a_n561_n139# a_303_73# a_n609_n42# a_n177_n139# a_n849_73# a_447_n42#
+ a_927_n42# a_n321_n42# a_879_73# a_n801_n42# a_159_n42# a_639_n42# a_n465_73# a_n513_n42#
+ a_n897_n42# a_783_n139# a_495_73# a_399_n139# a_351_n42# a_n33_n42# a_831_n42# a_n945_n139#
+ a_n225_n42# a_n705_n42# a_111_73# a_591_n139# a_543_n42# a_207_n139# a_n657_73#
+ VSUBS
X0 a_927_n42# a_879_73# a_831_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_73# a_n129_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_73# a_255_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_73# a_63_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n139# a_159_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_n139# a_351_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_543_n42# a_495_73# a_447_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_639_n42# a_591_n139# a_543_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_73# a_639_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n139# a_735_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n801_n42# a_n849_73# a_n897_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n513_n42# a_n561_n139# a_n609_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n321_n42# a_n369_n139# a_n417_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n225_n42# a_n273_73# a_n321_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n897_n42# a_n945_n139# a_n989_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X15 a_n705_n42# a_n753_n139# a_n801_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n609_n42# a_n657_73# a_n705_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n417_n42# a_n465_73# a_n513_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n139# a_n225_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_63_n42# a_15_n139# a_n33_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC45 a_63_n42# a_15_64# a_n417_n42# a_111_n130#
+ a_n273_n130# a_255_n42# a_n129_n42# a_n369_64# a_399_64# a_447_n42# a_n81_n130#
+ a_n321_n42# a_n509_n42# a_159_n42# a_351_n42# a_n33_n42# a_303_n130# a_n225_n42#
+ a_n177_64# a_207_64# a_n465_n130# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_n130# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_64# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n321_n42# a_n369_64# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n130# a_n509_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X8 a_n225_n42# a_n273_n130# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt buffer a_1504_1398# m5_n1320_776# a_n1158_1778# a_1504_1860# a_1596_1398#
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS w_1358_2156# m4_n1330_2222#
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552#
+ a_n1158_1778# a_n1158_1778# a_1436_1552# a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_n1158_1778# a_1436_1552# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_1436_1552# a_1436_1552# a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552#
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_n1158_1778# a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# a_n1158_1778#
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_1436_1552# a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1778# w_1358_2156# a_1436_1552# a_1436_1552#
+ w_1358_2156# a_1436_1552# a_n1158_1778# a_1436_1552# w_1358_2156# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ w_1358_2156# a_1436_1552# w_1358_2156# a_n1158_1778# w_1358_2156# w_1358_2156# w_1358_2156#
+ a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ a_1436_1552# w_1358_2156# a_n1158_1778# w_1358_2156# w_1358_2156# a_n1158_1778#
+ w_1358_2156# a_n1158_1778# w_1358_2156# a_1436_1552# a_1436_1552# a_1436_1552# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_1436_1552# w_1358_2156# w_1358_2156# a_n1158_1778#
+ a_n1158_1778# a_1436_1552# a_n1158_1778# a_1436_1552# a_1436_1552# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
X0 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X2 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X6 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X8 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X11 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X12 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X15 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X16 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X17 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X20 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X21 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X24 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X27 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X30 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X32 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X35 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X36 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X38 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X39 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X43 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X45 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X46 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X48 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X49 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X50 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X53 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
C0 a_1504_1860# a_1596_1398# 6.786759f
C1 a_1436_1552# a_1596_1398# 2.21286f
C2 a_1436_1552# w_1358_2156# 4.344402f
C3 a_1596_1398# a_1504_1398# 2.6505f
C4 m5_n1320_776# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 2.587544f
C5 a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 8.208134f
C6 w_1358_2156# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 6.120336f
C7 a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 9.825851f
.ends

.subckt sky130_fd_pr__pfet_01v8_X4L24Q a_n33_n126# w_n353_n226# a_n317_n126# a_n177_157#
+ a_159_n126# a_111_n223# a_n273_n223# a_255_n126# a_n129_n126# a_n81_n223# a_63_n126#
+ a_n225_n126# a_15_157# a_207_157# VSUBS
X0 a_159_n126# a_111_n223# a_63_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 a_n225_n126# a_n273_n223# a_n317_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X2 a_63_n126# a_15_157# a_n33_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 a_n129_n126# a_n177_157# a_n225_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_n33_n126# a_n81_n223# a_n129_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_255_n126# a_207_157# a_159_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_XJUN3E a_63_n42# a_15_64# a_111_n130# a_n273_n130#
+ a_255_n42# a_n129_n42# a_n317_n42# a_n81_n130# a_159_n42# a_n33_n42# a_n225_n42#
+ a_n177_64# a_207_64# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n225_n42# a_n273_n130# a_n317_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt and_gate a_514_134# w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206#
+ m1_748_n50#
Xsky130_fd_pr__pfet_01v8_X4L24Q_0 w_n260_286# w_n260_286# m1_748_n50# a_n78_396# w_n260_286#
+ a_n78_396# a_n78_396# m1_748_n50# m1_748_n50# a_n78_396# m1_748_n50# w_n260_286#
+ a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q
Xsky130_fd_pr__nfet_01v8_XJUN3E_0 m1_748_n50# a_n78_396# a_n78_396# a_n78_396# m1_748_n50#
+ m1_748_n50# m1_748_n50# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__nfet_01v8_XJUN3E
X0 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.1953 pd=1.57 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_n78_396# a_514_134# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X6 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 w_n260_286# a_514_134# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.1953 ps=1.57 w=1.26 l=0.15
X8 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X9 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X10 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X11 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 w_n260_286# a_n78_396# 3.023118f
C1 a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 2.455001f
C2 w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 6.963798f
.ends

.subckt buffer_and_gate in1 clk out gnd vdd
Xbuffer_0 gnd gnd clk vdd m1_5444_838# gnd vdd vdd buffer
Xand_gate_0 m1_5444_838# vdd gnd in1 out and_gate
C0 in1 gnd 2.619732f
C1 and_gate_0/a_n78_396# gnd 2.338147f
C2 clk gnd 8.795321f
C3 m1_5444_838# gnd 2.352718f
C4 vdd gnd 18.256077f
C5 buffer_0/a_1436_1552# gnd 11.512064f
.ends

.subckt capacito7 a_2858_n174# sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142# buffer_digital_0/i
+ a_5270_n124# m3_7758_166# buffer_and_gate_0/clk sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142#
+ m1_6370_n278# buffer_digital_0/VDD m1_602_n334# VSUBS
Xbuffer_digital_0 buffer_digital_0/i buffer_digital_0/in buffer_digital_0/VDD VSUBS
+ buffer_digital
Xsky130_fd_pr__pfet_01v8_4ZKXAA_0 m1_6370_n278# m1_6370_n278# VSUBS sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142#
+ m1_6370_n278# VSUBS m1_6370_n278# VSUBS m1_6370_n278# VSUBS VSUBS m1_6370_n278#
+ VSUBS m1_6370_n278# m1_6370_n278# VSUBS VSUBS m1_6370_n278# m1_6370_n278# VSUBS
+ m1_6370_n278# VSUBS VSUBS sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__nfet_01v8_9LGCGE_0 a_2858_n174# a_2858_n174# VSUBS VSUBS a_2858_n174#
+ VSUBS a_2858_n174# VSUBS a_2858_n174# VSUBS VSUBS VSUBS a_2858_n174# VSUBS VSUBS
+ a_2858_n174# VSUBS a_2858_n174# a_2858_n174# VSUBS a_2858_n174# a_2858_n174# VSUBS
+ VSUBS VSUBS VSUBS a_2858_n174# a_2858_n174# a_2858_n174# VSUBS a_2858_n174# a_2858_n174#
+ VSUBS VSUBS a_2858_n174# a_2858_n174# a_2858_n174# VSUBS VSUBS a_2858_n174# VSUBS
+ VSUBS sky130_fd_pr__nfet_01v8_9LGCGE
Xsky130_fd_pr__pfet_01v8_49FP49_0 m1_602_n334# m1_602_n334# VSUBS VSUBS m1_602_n334#
+ VSUBS sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142# m1_602_n334# m1_602_n334# VSUBS
+ VSUBS m1_602_n334# VSUBS VSUBS VSUBS m1_602_n334# VSUBS VSUBS m1_602_n334# m1_602_n334#
+ m1_602_n334# VSUBS m1_602_n334# m1_602_n334# m1_602_n334# VSUBS m1_602_n334# m1_602_n334#
+ VSUBS VSUBS VSUBS m1_602_n334# m1_602_n334# m1_602_n334# VSUBS m1_602_n334# m1_602_n334#
+ VSUBS VSUBS m1_602_n334# VSUBS VSUBS VSUBS sky130_fd_pr__pfet_01v8_49FP49
Xsky130_fd_pr__nfet_01v8_NJGC45_0 VSUBS a_5270_n124# VSUBS a_5270_n124# a_5270_n124#
+ VSUBS VSUBS a_5270_n124# a_5270_n124# VSUBS a_5270_n124# VSUBS VSUBS VSUBS VSUBS
+ VSUBS a_5270_n124# VSUBS a_5270_n124# a_5270_n124# a_5270_n124# VSUBS sky130_fd_pr__nfet_01v8_NJGC45
Xbuffer_and_gate_0 buffer_digital_0/in buffer_and_gate_0/clk buffer_and_gate_0/out
+ VSUBS buffer_digital_0/VDD buffer_and_gate
X0 buffer_and_gate_0/out m3_7758_166# sky130_fd_pr__cap_mim_m3_1 l=7.99 w=7.97
C0 buffer_digital_0/i buffer_digital_0/in 2.942645f
C1 m3_7758_166# VSUBS 2.50035f
C2 buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.473223f
C3 buffer_and_gate_0/clk VSUBS 8.924417f
C4 buffer_digital_0/VDD VSUBS 18.041912f
C5 buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.15507f
C6 a_5270_n124# VSUBS 3.420046f
C7 m1_602_n334# VSUBS 2.778242f
C8 a_2858_n174# VSUBS 6.69811f
C9 buffer_digital_0/in VSUBS 2.681842f
.ends

.subckt capacitor_8 capacitor_7_0/a_5270_n124# capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/clk
+ capacitor_7_0/buffer_digital_0/VDD capacitor_7_0/a_2858_n174# w_7118_n356# w_1380_n364#
+ VSUBS capacitor_7_0/buffer_digital_0/i
Xcapacitor_7_0 capacitor_7_0/a_2858_n174# w_7118_n356# capacitor_7_0/buffer_digital_0/i
+ capacitor_7_0/a_5270_n124# capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/clk
+ w_1380_n364# w_7118_n356# capacitor_7_0/buffer_digital_0/VDD w_1380_n364# VSUBS
+ capacito7
C0 capacitor_7_0/m3_7758_166# VSUBS 2.31534f
C1 capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C2 capacitor_7_0/buffer_and_gate_0/clk VSUBS 8.196827f
C3 capacitor_7_0/buffer_digital_0/VDD VSUBS 18.215277f
C4 capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C5 capacitor_7_0/a_5270_n124# VSUBS 2.356963f
C6 w_1380_n364# VSUBS 3.53509f
C7 capacitor_7_0/a_2858_n174# VSUBS 4.668162f
C8 capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
.ends

.subckt capacitors_1 clk1 capacitor_8_0/capacitor_7_0/a_2858_n174# capacitor_8_0/capacitor_7_0/a_5270_n124#
+ capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk capacitor_8_0/capacitor_7_0/buffer_digital_0/VDD
+ m1_7096_n308# capacitor_8_0/w_1380_n364# in1 VSUBS
Xcapacitor_8_0 capacitor_8_0/capacitor_7_0/a_5270_n124# clk1 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk
+ capacitor_8_0/capacitor_7_0/buffer_digital_0/VDD capacitor_8_0/capacitor_7_0/a_2858_n174#
+ m1_7096_n308# capacitor_8_0/w_1380_n364# VSUBS in1 capacitor_8
C0 clk1 VSUBS 2.376945f
C1 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C2 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk VSUBS 9.493001f
C3 capacitor_8_0/capacitor_7_0/buffer_digital_0/VDD VSUBS 22.92377f
C4 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C5 capacitor_8_0/capacitor_7_0/a_5270_n124# VSUBS 2.356963f
C6 capacitor_8_0/w_1380_n364# VSUBS 3.265198f
C7 capacitor_8_0/capacitor_7_0/a_2858_n174# VSUBS 4.668162f
C8 capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.613958f
.ends

.subckt sky130_fd_pr__pfet_01v8_4RPJ49 a_2031_73# a_1887_n42# a_3615_n42# a_3183_73#
+ a_n3729_73# a_n2529_n42# a_1503_n42# a_63_n42# a_n753_n139# a_n3393_n42# a_n369_n139#
+ a_n1425_73# a_n1281_n42# a_n2961_73# a_687_73# a_n2577_73# a_n417_n42# a_2367_n42#
+ a_n1761_n42# a_n3009_n42# a_n2673_n139# a_2847_n42# a_n2289_n139# a_n3633_n139#
+ a_2607_73# a_n3249_n139# a_n1713_n139# a_3759_73# a_n1329_n139# a_255_n42# a_1455_73#
+ a_n2241_n42# a_2991_73# a_3471_n139# a_735_n42# a_1551_n139# a_3087_n139# a_1599_n42#
+ a_3327_n42# a_1167_n139# a_n2721_n42# a_n81_73# a_2511_n139# a_1215_n42# a_n273_73#
+ a_2127_n139# a_n993_n42# a_3807_n42# a_15_n139# a_303_73# a_n3585_n42# a_n129_n42#
+ a_2079_n42# a_n561_n139# a_n3345_73# a_n3201_n42# a_n1473_n42# a_n177_n139# a_n1041_73#
+ a_n609_n42# a_2559_n42# a_n2193_73# a_n1953_n42# a_n849_73# w_n3905_n142# a_n2481_n139#
+ a_n2097_n139# a_n3441_n139# a_1791_n42# a_n1521_n139# a_n3057_n139# a_2223_73# a_447_n42#
+ a_3039_n42# a_n1137_n139# a_3375_73# a_n2433_n42# a_927_n42# a_1071_73# a_n1617_73#
+ a_n2913_n42# a_3519_n42# a_975_n139# a_879_73# a_n2769_73# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n1185_n42# a_n801_n42# a_n3777_n42# a_2751_n42# a_n1665_n42#
+ a_1647_73# a_2799_73# a_3231_n42# a_159_n42# a_n2145_n42# a_n465_73# a_1983_n42#
+ a_3711_n42# a_639_n42# a_n2625_n42# a_1119_n42# a_n3537_73# a_n897_n42# a_n513_n42#
+ a_n1233_73# a_n3489_n42# a_2463_n42# a_783_n139# a_495_73# a_399_n139# a_n2385_73#
+ a_2895_n139# a_n3105_n42# a_n1377_n42# a_2943_n42# a_1935_n139# a_n1857_n42# a_351_n42#
+ a_2415_73# a_n33_n42# a_3567_73# a_831_n42# a_1695_n42# a_3423_n42# a_1263_73# a_n945_n139#
+ a_n2337_n42# a_1311_n42# a_n1809_73# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2175_n42#
+ a_n2865_n139# a_n1089_n42# a_n3825_n139# a_111_73# a_n2001_73# a_n3869_n42# a_n705_n42#
+ a_2655_n42# a_n1905_n139# a_n3153_73# a_591_n139# a_1839_73# a_n1569_n42# a_3663_n139#
+ a_1743_n139# a_3279_n139# a_543_n42# a_207_n139# a_n657_73# a_1359_n139# a_2703_n139#
+ a_3135_n42# VSUBS a_2319_n139# a_n2049_n42# a_1023_n42#
X0 a_n2241_n42# a_n2289_n139# a_n2337_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n2913_n42# a_n2961_73# a_n3009_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n2721_n42# a_n2769_73# a_n2817_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n2625_n42# a_n2673_n139# a_n2721_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n2433_n42# a_n2481_n139# a_n2529_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n2337_n42# a_n2385_73# a_n2433_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n2145_n42# a_n2193_73# a_n2241_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n2049_n42# a_n2097_n139# a_n2145_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n2817_n42# a_n2865_n139# a_n2913_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n2529_n42# a_n2577_73# a_n2625_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_2079_n42# a_2031_73# a_1983_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_2175_n42# a_2127_n139# a_2079_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_2271_n42# a_2223_73# a_2175_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_2367_n42# a_2319_n139# a_2271_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_2463_n42# a_2415_73# a_2367_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_2655_n42# a_2607_73# a_2559_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_2751_n42# a_2703_n139# a_2655_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_2943_n42# a_2895_n139# a_2847_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_2559_n42# a_2511_n139# a_2463_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_2847_n42# a_2799_73# a_2751_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_927_n42# a_879_73# a_831_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_1023_n42# a_975_n139# a_927_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n1953_n42# a_n2001_73# a_n2049_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_n1761_n42# a_n1809_73# a_n1857_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n1665_n42# a_n1713_n139# a_n1761_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n1857_n42# a_n1905_n139# a_n1953_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n1569_n42# a_n1617_73# a_n1665_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_1119_n42# a_1071_73# a_1023_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1215_n42# a_1167_n139# a_1119_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1311_n42# a_1263_73# a_1215_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_1407_n42# a_1359_n139# a_1311_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1503_n42# a_1455_73# a_1407_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_1695_n42# a_1647_73# a_1599_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1791_n42# a_1743_n139# a_1695_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1599_n42# a_1551_n139# a_1503_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_1887_n42# a_1839_73# a_1791_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_1983_n42# a_1935_n139# a_1887_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n33_n42# a_n81_73# a_n129_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_351_n42# a_303_73# a_255_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_159_n42# a_111_73# a_63_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_255_n42# a_207_n139# a_159_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_447_n42# a_399_n139# a_351_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_543_n42# a_495_73# a_447_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_639_n42# a_591_n139# a_543_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_735_n42# a_687_73# a_639_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_831_n42# a_783_n139# a_735_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_n1473_n42# a_n1521_n139# a_n1569_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_n1377_n42# a_n1425_73# a_n1473_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_n1281_n42# a_n1329_n139# a_n1377_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_n1185_n42# a_n1233_73# a_n1281_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n1089_n42# a_n1137_n139# a_n1185_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_n993_n42# a_n1041_73# a_n1089_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_n801_n42# a_n849_73# a_n897_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_n513_n42# a_n561_n139# a_n609_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_n321_n42# a_n369_n139# a_n417_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_n225_n42# a_n273_73# a_n321_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_n897_n42# a_n945_n139# a_n993_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_n705_n42# a_n753_n139# a_n801_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_n609_n42# a_n657_73# a_n705_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n417_n42# a_n465_73# a_n513_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n129_n42# a_n177_n139# a_n225_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_3327_n42# a_3279_n139# a_3231_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_3423_n42# a_3375_73# a_3327_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_3615_n42# a_3567_73# a_3519_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_3711_n42# a_3663_n139# a_3615_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_3519_n42# a_3471_n139# a_3423_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_3807_n42# a_3759_73# a_3711_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n3201_n42# a_n3249_n139# a_n3297_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_63_n42# a_15_n139# a_n33_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n3681_n42# a_n3729_73# a_n3777_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n3585_n42# a_n3633_n139# a_n3681_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n3393_n42# a_n3441_n139# a_n3489_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n3297_n42# a_n3345_73# a_n3393_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n3105_n42# a_n3153_73# a_n3201_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_n3009_n42# a_n3057_n139# a_n3105_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3231_n42# a_3183_73# a_3135_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_n3777_n42# a_n3825_n139# a_n3869_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X77 a_n3489_n42# a_n3537_73# a_n3585_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3039_n42# a_2991_73# a_2943_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3135_n42# a_3087_n139# a_3039_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 w_n3905_n142# VSUBS 6.63223f
.ends

.subckt sky130_fd_pr__pfet_01v8_E9H44Q a_15_n42# a_n15_n68# w_n109_n104# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# w_n109_n104# sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_9AYYDL a_n158_n300# w_n194_n362# a_100_n300# a_n100_n326#
+ VSUBS
X0 a_100_n300# a_n100_n326# a_n158_n300# w_n194_n362# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt pmos_cp1 a_168_22# m1_532_58# w_n14_n142# a_424_18# m1_14_56# VSUBS
Xsky130_fd_pr__pfet_01v8_E9H44Q_0 w_n14_n142# a_168_22# w_n14_n142# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_E9H44Q_1 a_168_22# a_424_18# w_n14_n142# w_n14_n142# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_9AYYDL_0 m1_14_56# w_n14_n142# w_n14_n142# a_168_22# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
Xsky130_fd_pr__pfet_01v8_9AYYDL_1 w_n14_n142# w_n14_n142# m1_532_58# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
C0 w_n14_n142# VSUBS 2.470929f
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC8F a_15_n130# a_1887_n42# a_3615_n42# a_1647_64#
+ a_n561_n130# a_n2529_n42# a_1503_n42# a_2799_64# a_63_n42# a_n177_n130# a_n3393_n42#
+ a_n1281_n42# a_n465_64# a_n417_n42# a_2367_n42# a_n1761_n42# a_n2481_n130# a_n3009_n42#
+ a_n2097_n130# a_n3441_n130# a_2847_n42# a_n1521_n130# a_n3057_n130# a_n3537_64#
+ a_n1137_n130# a_255_n42# a_n1233_64# a_495_64# a_n2241_n42# a_n2385_64# a_975_n130#
+ a_735_n42# a_1599_n42# a_3327_n42# a_n2721_n42# a_1215_n42# a_2415_64# a_n993_n42#
+ a_3807_n42# a_3567_64# a_n3585_n42# a_n129_n42# a_2079_n42# a_1263_64# a_n3201_n42#
+ a_n1473_n42# a_n1809_64# a_n609_n42# a_2559_n42# a_n1953_n42# a_111_64# a_n2001_64#
+ a_1791_n42# a_447_n42# a_n3153_64# a_3039_n42# a_n2433_n42# a_1839_64# a_927_n42#
+ a_n2913_n42# a_3519_n42# a_783_n130# a_399_n130# a_2895_n130# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n657_64# a_n1185_n42# a_1935_n130# a_n801_n42# a_2031_64#
+ a_n3777_n42# a_2751_n42# a_3183_64# a_n1665_n42# a_n3729_64# a_n1425_64# a_687_64#
+ a_n2961_64# a_n945_n130# a_n2577_64# a_3231_n42# a_159_n42# a_n2145_n42# a_1983_n42#
+ a_3711_n42# a_2607_64# a_639_n42# a_n2625_n42# a_3759_64# a_n2865_n130# a_1119_n42#
+ a_n3825_n130# a_1455_64# a_n1905_n130# a_2991_64# a_n897_n42# a_591_n130# a_n513_n42#
+ a_n3489_n42# a_2463_n42# a_n3105_n42# a_n1377_n42# a_n81_64# a_n273_64# a_3663_n130#
+ a_3279_n130# a_2943_n42# a_1743_n130# a_207_n130# a_2703_n130# a_1359_n130# a_n1857_n42#
+ a_2319_n130# a_351_n42# a_303_64# a_n3345_64# a_n33_n42# a_831_n42# a_n1041_64#
+ a_1695_n42# a_3423_n42# a_n753_n130# a_n369_n130# a_n2193_64# a_n2337_n42# a_1311_n42#
+ a_n849_64# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2223_64# a_n2673_n130# a_2175_n42#
+ a_3375_64# a_n2289_n130# a_n3633_n130# a_n1089_n42# a_n3249_n130# a_n1713_n130#
+ a_n3869_n42# a_n705_n42# a_2655_n42# a_1071_64# a_n1329_n130# a_n1617_64# a_n1569_n42#
+ a_879_64# a_n2769_64# a_3471_n130# a_3087_n130# a_1551_n130# a_2511_n130# a_543_n42#
+ a_1167_n130# a_3135_n42# a_2127_n130# VSUBS a_n2049_n42# a_1023_n42#
X0 a_n3201_n42# a_n3249_n130# a_n3297_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n3681_n42# a_n3729_64# a_n3777_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n3585_n42# a_n3633_n130# a_n3681_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n3393_n42# a_n3441_n130# a_n3489_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n3297_n42# a_n3345_64# a_n3393_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n3105_n42# a_n3153_64# a_n3201_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n3009_n42# a_n3057_n130# a_n3105_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n3777_n42# a_n3825_n130# a_n3869_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X9 a_n3489_n42# a_n3537_64# a_n3585_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_3135_n42# a_3087_n130# a_3039_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_3231_n42# a_3183_64# a_3135_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_3039_n42# a_2991_64# a_2943_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n2241_n42# a_n2289_n130# a_n2337_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n2913_n42# a_n2961_64# a_n3009_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n2721_n42# a_n2769_64# a_n2817_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n2625_n42# a_n2673_n130# a_n2721_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n2433_n42# a_n2481_n130# a_n2529_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n2337_n42# a_n2385_64# a_n2433_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n2145_n42# a_n2193_64# a_n2241_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_n2049_n42# a_n2097_n130# a_n2145_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n2817_n42# a_n2865_n130# a_n2913_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n2529_n42# a_n2577_64# a_n2625_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2175_n42# a_2127_n130# a_2079_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_2271_n42# a_2223_64# a_2175_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2463_n42# a_2415_64# a_2367_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_2751_n42# a_2703_n130# a_2655_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_2079_n42# a_2031_64# a_1983_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_2367_n42# a_2319_n130# a_2271_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2559_n42# a_2511_n130# a_2463_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_2655_n42# a_2607_64# a_2559_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_2847_n42# a_2799_64# a_2751_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_2943_n42# a_2895_n130# a_2847_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1023_n42# a_975_n130# a_927_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_n1953_n42# a_n2001_64# a_n2049_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_n1761_n42# a_n1809_64# a_n1857_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n1665_n42# a_n1713_n130# a_n1761_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_n1857_n42# a_n1905_n130# a_n1953_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_n1569_n42# a_n1617_64# a_n1665_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1215_n42# a_1167_n130# a_1119_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1311_n42# a_1263_64# a_1215_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1503_n42# a_1455_64# a_1407_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_1791_n42# a_1743_n130# a_1695_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1119_n42# a_1071_64# a_1023_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_1407_n42# a_1359_n130# a_1311_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_1599_n42# a_1551_n130# a_1503_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1695_n42# a_1647_64# a_1599_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_1887_n42# a_1839_64# a_1791_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_1983_n42# a_1935_n130# a_1887_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n1473_n42# a_n1521_n130# a_n1569_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n1281_n42# a_n1329_n130# a_n1377_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_n1185_n42# a_n1233_64# a_n1281_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_n993_n42# a_n1041_64# a_n1089_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_n1377_n42# a_n1425_64# a_n1473_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_n1089_n42# a_n1137_n130# a_n1185_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n897_n42# a_n945_n130# a_n993_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_3327_n42# a_3279_n130# a_3231_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3423_n42# a_3375_64# a_3327_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_3615_n42# a_3567_64# a_3519_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X77 a_3711_n42# a_3663_n130# a_3615_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3519_n42# a_3471_n130# a_3423_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3807_n42# a_3759_64# a_3711_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt charge_pump1 clk_in input1 input2 in1 in2 in6 in7 g1 g2 clk clkb m1_12464_n576#
+ a_3340_18086# in4 in3 in5 in8 vin vdd gnd
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 g1 clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 g2 clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 vin input1 input2 g1 g2 vin gnd nmos_dnw3
Xclock_0 clk_in vdd gnd clk clkb clock
Xcapacitor_8_0 vdd input1 clk vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 clkb vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 vdd vdd clk vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_1 input2 vdd vdd clkb vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_2 input1 vdd vdd clk vdd vdd vdd in2 gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 vdd vdd clk vdd vdd vdd in3 gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_4 input2 vdd vdd clkb vdd vdd vdd in2 gnd capacitors_1
Xcapacitors_1_5 input2 vdd vdd clkb vdd vdd vdd in3 gnd capacitors_1
Xcapacitors_1_6 input1 vdd vdd clk vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_7 input1 vdd vdd clk vdd vdd vdd in5 gnd capacitors_1
Xcapacitors_1_8 input1 vdd vdd clk vdd vdd vdd in6 gnd capacitors_1
Xcapacitors_1_9 input1 vdd vdd clk vdd vdd vdd in7 gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 vdd vdd clkb vdd vdd vdd in7 gnd capacitors_1
Xcapacitors_1_11 input2 vdd vdd clkb vdd vdd vdd in6 gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 vdd vdd clkb vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_12 input2 vdd vdd clkb vdd vdd vdd in5 gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clkb input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clk input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 clk m1_12464_n576# 2.312213f
C1 vdd clkb 26.212053f
C2 input2 input1 3.059187f
C3 vdd input1 26.823656f
C4 vdd clk 32.205326f
C5 vin vdd 9.1372f
C6 vin clk 2.188878f
C7 vdd input2 26.500195f
C8 clkb m1_12464_n576# 2.207061f
C9 input1 gnd 30.964584f
C10 input2 gnd 31.05456f
C11 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.396566f
C12 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.07966f
C13 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634299f
C14 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398093f
C15 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.08029f
C16 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633591f
C17 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.392522f
C18 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079402f
C19 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634253f
C20 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398324f
C21 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079739f
C22 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633955f
C23 m1_4341_n519# gnd 4.097057f
C24 m1_12659_300# gnd 2.789905f
C25 m1_12464_n576# gnd 5.227879f
C26 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.397358f
C27 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079556f
C28 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634405f
C29 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.394424f
C30 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079654f
C31 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634067f
C32 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393486f
C33 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.07973f
C34 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633915f
C35 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393389f
C36 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079822f
C37 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633871f
C38 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398049f
C39 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079473f
C40 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633938f
C41 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.396035f
C42 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079795f
C43 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634021f
C44 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.395022f
C45 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079731f
C46 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634052f
C47 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.392135f
C48 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.078752f
C49 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633513f
C50 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.338151f
C51 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.97841f
C52 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61055f
C53 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.33782f
C54 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978384f
C55 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.610197f
C56 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393725f
C57 clkb gnd 91.86899f
C58 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.080707f
C59 capacitor_8_1/capacitor_7_0/buffer_digital_0/in gnd 2.639488f
C60 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.397516f
C61 clk gnd 91.63095f
C62 vdd gnd 0.653035p
C63 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079217f
C64 capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.639593f
C65 clock_0/a_2432_n962# gnd 8.68424f **FLOATING
C66 clock_0/a_2020_n482# gnd 2.567662f **FLOATING
C67 clock_0/a_344_102# gnd 2.813001f
C68 clock_0/a_2402_572# gnd 2.172722f
C69 clock_0/a_344_n986# gnd 2.381627f
C70 clock_0/a_3246_118# gnd 6.834443f
C71 g2 gnd 2.344427f
C72 vin gnd 10.416249f
.ends

.subckt sky130_fd_pr__nfet_01v8_TKGCLY a_n1425_n130# a_1887_n42# a_1503_n42# a_63_n42#
+ a_15_64# a_2127_64# a_n1281_n42# a_111_n130# a_879_n130# a_1263_n130# a_n417_n42#
+ a_2367_n42# a_2223_n130# a_n1761_n42# a_n1905_64# a_n273_n130# a_255_n42# a_n2241_n42#
+ a_735_n42# a_1599_n42# a_1935_64# a_n2429_n42# a_1215_n42# a_n2193_n130# a_n993_n42#
+ a_n1233_n130# a_n753_64# a_n369_64# a_n129_n42# a_2079_n42# a_n1473_n42# a_n609_n42#
+ a_687_n130# a_1071_n130# a_n1953_n42# a_2031_n130# a_n1521_64# a_n1137_64# a_783_64#
+ a_399_64# a_1839_n130# a_n2289_64# a_1791_n42# a_447_n42# a_927_n42# a_n81_n130#
+ a_2319_64# a_n849_n130# a_n321_n42# a_1407_n42# a_1551_64# a_2271_n42# a_1167_64#
+ a_n1185_n42# a_n801_n42# a_n1041_n130# a_n2001_n130# a_n1665_n42# a_n1809_n130#
+ a_495_n130# a_159_n42# a_n2145_n42# a_1647_n130# a_1983_n42# a_639_n42# a_n945_64#
+ a_1119_n42# a_n897_n42# a_n657_n130# a_n513_n42# a_n1377_n42# a_n1713_64# a_n1329_64#
+ a_975_64# a_n1857_n42# a_351_n42# a_n33_n42# a_n1617_n130# a_831_n42# a_1695_n42#
+ a_n2337_n42# a_1311_n42# a_303_n130# a_1743_64# a_1359_64# a_1455_n130# a_n225_n42#
+ a_2175_n42# a_n561_64# a_n1089_n42# a_n177_64# a_n705_n42# a_n465_n130# a_n1569_n42#
+ a_207_64# a_543_n42# a_591_64# a_n2097_64# a_n2385_n130# VSUBS a_n2049_n42# a_1023_n42#
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n2241_n42# a_n2289_64# a_n2337_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n2337_n42# a_n2385_n130# a_n2429_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3 a_n2145_n42# a_n2193_n130# a_n2241_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n2049_n42# a_n2097_64# a_n2145_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_2175_n42# a_2127_64# a_2079_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_2271_n42# a_2223_n130# a_2175_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_2079_n42# a_2031_n130# a_1983_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_2367_n42# a_2319_64# a_2271_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_927_n42# a_879_n130# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_1023_n42# a_975_64# a_927_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n1953_n42# a_n2001_n130# a_n2049_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n1761_n42# a_n1809_n130# a_n1857_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n1665_n42# a_n1713_64# a_n1761_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n1857_n42# a_n1905_64# a_n1953_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n1569_n42# a_n1617_n130# a_n1665_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_1215_n42# a_1167_64# a_1119_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_1311_n42# a_1263_n130# a_1215_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_1503_n42# a_1455_n130# a_1407_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_1791_n42# a_1743_64# a_1695_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_1119_n42# a_1071_n130# a_1023_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_1407_n42# a_1359_64# a_1311_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1599_n42# a_1551_64# a_1503_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_1695_n42# a_1647_n130# a_1599_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_1887_n42# a_1839_n130# a_1791_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_1983_n42# a_1935_64# a_1887_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_351_n42# a_303_n130# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_447_n42# a_399_64# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_543_n42# a_495_n130# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_735_n42# a_687_n130# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_831_n42# a_783_64# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_639_n42# a_591_64# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_n1473_n42# a_n1521_64# a_n1569_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_n1281_n42# a_n1329_64# a_n1377_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n1185_n42# a_n1233_n130# a_n1281_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_n993_n42# a_n1041_n130# a_n1089_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_n1377_n42# a_n1425_n130# a_n1473_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_n1089_n42# a_n1137_64# a_n1185_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_n321_n42# a_n369_64# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_n801_n42# a_n849_n130# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_n705_n42# a_n753_64# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_n609_n42# a_n657_n130# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_n513_n42# a_n561_64# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_n417_n42# a_n465_n130# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_n225_n42# a_n273_n130# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_n897_n42# a_n945_64# a_n993_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt nmos_decap_10 a_n2_210# m1_n10_n42# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGC45_0 m1_n10_n42# a_n2_210# m1_n10_n42# a_n2_210# a_n2_210#
+ m1_n10_n42# m1_n10_n42# a_n2_210# a_n2_210# m1_n10_n42# a_n2_210# m1_n10_n42# m1_n10_n42#
+ m1_n10_n42# m1_n10_n42# m1_n10_n42# a_n2_210# m1_n10_n42# a_n2_210# a_n2_210# a_n2_210#
+ VSUBS sky130_fd_pr__nfet_01v8_NJGC45
C0 a_n2_210# VSUBS 2.327241f
.ends

.subckt pmos_decap_10 a_12_230# w_6_4# VSUBS
Xsky130_fd_pr__pfet_01v8_4ZKXAA_0 w_6_4# w_6_4# a_12_230# w_6_4# w_6_4# a_12_230#
+ w_6_4# a_12_230# w_6_4# a_12_230# a_12_230# w_6_4# a_12_230# w_6_4# w_6_4# a_12_230#
+ a_12_230# w_6_4# w_6_4# a_12_230# w_6_4# a_12_230# VSUBS sky130_fd_pr__pfet_01v8_4ZKXAA
.ends

.subckt cp1_buffer1 charge_pump1_0/in8 charge_pump1_0/in4 charge_pump1_0/in3 charge_pump1_0/in5
+ charge_pump1_0/in2 charge_pump1_0/vin charge_pump1_0/in6 clk_out clk_in charge_pump1_0/in1
+ charge_pump1_0/m1_12464_n576# charge_pump1_0/in7 gnd vdd
Xsky130_fd_pr__nfet_01v8_HRDN5X_0 vdd gnd vdd vdd vdd vdd gnd gnd gnd vdd gnd vdd
+ gnd gnd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd gnd gnd gnd gnd vdd gnd
+ sky130_fd_pr__nfet_01v8_HRDN5X
Xcharge_pump1_0 clk_out charge_pump1_0/input1 charge_pump1_0/input2 charge_pump1_0/in1
+ charge_pump1_0/in2 charge_pump1_0/in6 charge_pump1_0/in7 charge_pump1_0/g1 charge_pump1_0/g2
+ charge_pump1_0/clk charge_pump1_0/clkb charge_pump1_0/m1_12464_n576# gnd charge_pump1_0/in4
+ charge_pump1_0/in3 charge_pump1_0/in5 charge_pump1_0/in8 charge_pump1_0/vin vdd
+ gnd charge_pump1
Xsky130_fd_pr__nfet_01v8_TKGCLY_0 vdd gnd gnd gnd vdd vdd gnd vdd vdd vdd gnd gnd
+ vdd gnd vdd vdd gnd gnd gnd gnd vdd gnd gnd vdd gnd vdd vdd vdd gnd gnd gnd gnd
+ vdd vdd gnd vdd vdd vdd vdd vdd vdd vdd gnd gnd gnd vdd vdd vdd gnd gnd vdd gnd
+ vdd gnd gnd vdd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd gnd gnd vdd gnd gnd vdd
+ vdd vdd gnd gnd gnd vdd gnd gnd gnd gnd vdd vdd vdd vdd gnd gnd vdd gnd vdd gnd
+ vdd gnd vdd gnd vdd vdd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_TKGCLY
Xbuffer_digital_0 clk_int clk_out vdd gnd buffer_digital
Xbuffer_digital_1 clk_in clk_int vdd gnd buffer_digital
Xnmos_decap_10_0 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_1 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_2 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_3 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_4 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_6 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_5 vdd gnd gnd nmos_decap_10
Xpmos_decap_10_0 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_1 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_2 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_3 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_4 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_5 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_6 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_7 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_9 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_8 gnd vdd gnd pmos_decap_10
C0 vdd clk_out 5.285868f
C1 clk_in gnd 6.708698f
C2 clk_out gnd 13.128814f
C3 charge_pump1_0/input1 gnd 22.463037f
C4 charge_pump1_0/input2 gnd 22.175129f
C5 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C6 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C7 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C8 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C9 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C10 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C11 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C12 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C13 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C14 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C15 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C16 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C17 charge_pump1_0/m1_4341_n519# gnd 3.771611f
C18 charge_pump1_0/m1_12659_300# gnd 2.538747f
C19 charge_pump1_0/m1_12464_n576# gnd 4.33476f
C20 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C21 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C22 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C23 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C24 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C25 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C26 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C27 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C28 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C29 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C30 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C31 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C32 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C33 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C34 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C35 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C36 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C37 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C38 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C39 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C40 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C41 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C42 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C43 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C44 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C45 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C46 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C47 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C48 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C49 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C50 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C51 charge_pump1_0/clkb gnd 90.01183f
C52 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C53 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C54 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.337696f
C55 charge_pump1_0/clk gnd 89.583115f
C56 vdd gnd 0.575054p
C57 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978376f
C58 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.608221f
C59 charge_pump1_0/clock_0/a_2432_n962# gnd 8.68424f **FLOATING
C60 charge_pump1_0/clock_0/a_2020_n482# gnd 2.56615f **FLOATING
C61 charge_pump1_0/clock_0/a_344_102# gnd 2.809951f
C62 charge_pump1_0/clock_0/a_2402_572# gnd 2.172722f
C63 charge_pump1_0/clock_0/a_344_n986# gnd 2.381627f
C64 charge_pump1_0/clock_0/a_3246_118# gnd 6.834443f
C65 charge_pump1_0/g2 gnd 2.344427f
C66 charge_pump1_0/vin gnd 10.376139f
.ends

.subckt charge_pump1_reverse input1 input2 in1 in2 in6 in7 vdd m1_12464_n576# clock_1/clk_in
+ a_3340_18086# in4 in3 in5 gnd in8 nmos_dnw3_0/vs
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 nmos_dnw3_0/vs input1 input2 nmos_dnw3_0/clk nmos_dnw3_0/clkb nmos_dnw3_0/vs
+ gnd nmos_dnw3
Xclock_1 clock_1/clk_in vdd gnd clock_1/clk clock_1/clkb clock
Xcapacitor_8_0 vdd input1 clock_1/clkb vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 clock_1/clk vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 vdd vdd clock_1/clkb vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_1 input2 vdd vdd clock_1/clk vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_2 input1 vdd vdd clock_1/clkb vdd vdd vdd in2 gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 vdd vdd clock_1/clkb vdd vdd vdd in3 gnd capacitors_1
Xcapacitors_1_4 input2 vdd vdd clock_1/clk vdd vdd vdd in2 gnd capacitors_1
Xcapacitors_1_5 input2 vdd vdd clock_1/clk vdd vdd vdd in3 gnd capacitors_1
Xcapacitors_1_6 input1 vdd vdd clock_1/clkb vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_7 input1 vdd vdd clock_1/clkb vdd vdd vdd in5 gnd capacitors_1
Xcapacitors_1_8 input1 vdd vdd clock_1/clkb vdd vdd vdd in6 gnd capacitors_1
Xcapacitors_1_9 input1 vdd vdd clock_1/clkb vdd vdd vdd in7 gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 vdd vdd clock_1/clk vdd vdd vdd in7 gnd capacitors_1
Xcapacitors_1_11 input2 vdd vdd clock_1/clk vdd vdd vdd in6 gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 vdd vdd clock_1/clk vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_12 input2 vdd vdd clock_1/clk vdd vdd vdd in5 gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clock_1/clk input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clock_1/clkb input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 vdd clock_1/clk 28.684513f
C1 input2 input1 3.059187f
C2 input1 vdd 26.538095f
C3 nmos_dnw3_0/vs clock_1/clkb 2.218511f
C4 m1_12464_n576# clock_1/clk 2.140857f
C5 nmos_dnw3_0/vs vdd 9.238383f
C6 vdd clock_1/clkb 32.26193f
C7 input2 vdd 26.544638f
C8 m1_12464_n576# clock_1/clkb 2.29778f
C9 input1 gnd 31.198782f
C10 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.396567f
C11 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079662f
C12 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634299f
C13 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398093f
C14 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.080289f
C15 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633591f
C16 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.392522f
C17 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079402f
C18 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634253f
C19 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398324f
C20 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079739f
C21 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633955f
C22 m1_4341_n519# gnd 3.765437f
C23 input2 gnd 30.578617f
C24 m1_12659_300# gnd 3.025714f
C25 m1_12464_n576# gnd 5.503336f
C26 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.397358f
C27 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079556f
C28 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634405f
C29 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.394424f
C30 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079656f
C31 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634067f
C32 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393486f
C33 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079731f
C34 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633915f
C35 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39339f
C36 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.07982f
C37 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633871f
C38 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398049f
C39 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079472f
C40 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633938f
C41 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.396035f
C42 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079795f
C43 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634021f
C44 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.395022f
C45 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079731f
C46 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634052f
C47 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.392135f
C48 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.078753f
C49 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633513f
C50 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.338151f
C51 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.97841f
C52 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61055f
C53 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.33782f
C54 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978384f
C55 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.610197f
C56 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393725f
C57 clock_1/clk gnd 96.75779f
C58 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.080708f
C59 capacitor_8_1/capacitor_7_0/buffer_digital_0/in gnd 2.639487f
C60 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.397516f
C61 clock_1/clkb gnd 0.104535p
C62 vdd gnd 0.659544p
C63 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079217f
C64 capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.639594f
C65 clock_1/a_2432_n962# gnd 8.693805f **FLOATING
C66 clock_1/a_2020_n482# gnd 2.56615f **FLOATING
C67 clock_1/a_344_102# gnd 2.809951f
C68 clock_1/a_2402_572# gnd 2.172722f
C69 clock_1/a_344_n986# gnd 2.381627f
C70 clock_1/a_3246_118# gnd 6.834443f
C71 nmos_dnw3_0/vs gnd 10.39343f
.ends

.subckt cp1_buffer1_reverse charge_pump1_reverse_0/m1_12464_n576# charge_pump1_reverse_0/in6
+ charge_pump1_reverse_0/in7 charge_pump1_reverse_0/in1 buffer_digital_0/in charge_pump1_reverse_0/in8
+ buffer_digital_1/VDD charge_pump1_reverse_0/nmos_dnw3_0/vs charge_pump1_reverse_0/in4
+ charge_pump1_reverse_0/in3 buffer_digital_1/i charge_pump1_reverse_0/in5 charge_pump1_reverse_0/in2
+ VSUBS
Xpmos_decap_10_10 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_11 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_12 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_13 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_14 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xcharge_pump1_reverse_0 charge_pump1_reverse_0/input1 charge_pump1_reverse_0/input2
+ charge_pump1_reverse_0/in1 charge_pump1_reverse_0/in2 charge_pump1_reverse_0/in6
+ charge_pump1_reverse_0/in7 buffer_digital_1/VDD charge_pump1_reverse_0/m1_12464_n576#
+ buffer_digital_0/in VSUBS charge_pump1_reverse_0/in4 charge_pump1_reverse_0/in3
+ charge_pump1_reverse_0/in5 VSUBS charge_pump1_reverse_0/in8 charge_pump1_reverse_0/nmos_dnw3_0/vs
+ charge_pump1_reverse
Xbuffer_digital_0 buffer_digital_0/i buffer_digital_0/in buffer_digital_1/VDD VSUBS
+ buffer_digital
Xbuffer_digital_1 buffer_digital_1/i buffer_digital_0/i buffer_digital_1/VDD VSUBS
+ buffer_digital
Xnmos_decap_10_0 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_1 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_2 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_3 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_4 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_10 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_11 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_5 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_6 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_12 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_7 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_8 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_0 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xnmos_decap_10_9 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_1 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_2 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_3 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_4 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_5 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_6 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_7 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_9 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_8 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
C0 buffer_digital_1/VDD buffer_digital_0/in 5.980218f
C1 buffer_digital_1/VDD charge_pump1_reverse_0/clock_1/clkb 2.735452f
C2 buffer_digital_1/i VSUBS 6.664738f
C3 charge_pump1_reverse_0/input1 VSUBS 22.596436f
C4 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C5 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C6 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C7 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C8 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C9 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C10 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C11 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C12 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C13 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C14 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C15 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C16 charge_pump1_reverse_0/m1_4341_n519# VSUBS 3.33176f
C17 charge_pump1_reverse_0/input2 VSUBS 22.21436f
C18 charge_pump1_reverse_0/m1_12659_300# VSUBS 2.683598f
C19 charge_pump1_reverse_0/m1_12464_n576# VSUBS 4.637158f
C20 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C21 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C22 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C23 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C24 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C25 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C26 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C27 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C28 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C29 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C30 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C31 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C32 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C33 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C34 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C35 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C36 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C37 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C38 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C39 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C40 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C41 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C42 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C43 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C44 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C45 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C46 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C47 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C48 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C49 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C50 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C51 charge_pump1_reverse_0/clock_1/clk VSUBS 94.69408f
C52 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C53 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C54 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C55 charge_pump1_reverse_0/clock_1/clkb VSUBS 0.101101p
C56 buffer_digital_1/VDD VSUBS 0.574874p
C57 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C58 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C59 charge_pump1_reverse_0/clock_1/a_2432_n962# VSUBS 8.68424f **FLOATING
C60 charge_pump1_reverse_0/clock_1/a_2020_n482# VSUBS 2.56615f **FLOATING
C61 charge_pump1_reverse_0/clock_1/a_344_102# VSUBS 2.809951f
C62 charge_pump1_reverse_0/clock_1/a_2402_572# VSUBS 2.172722f
C63 charge_pump1_reverse_0/clock_1/a_344_n986# VSUBS 2.381632f
C64 buffer_digital_0/in VSUBS 16.517464f
C65 charge_pump1_reverse_0/clock_1/a_3246_118# VSUBS 6.834443f
C66 charge_pump1_reverse_0/nmos_dnw3_0/vs VSUBS 10.345203f
.ends

.subckt cp1_buffer_5stage cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/in8
+ cp1_buffer1_2/charge_pump1_0/in7 cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/m1_12464_n576# cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_0/clk_in cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_0/charge_pump1_0/vin cp1_buffer1_1/charge_pump1_0/vin cp1_buffer1_2/vdd
+ VSUBS cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/vin
Xcp1_buffer1_0 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_0/charge_pump1_0/vin
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_0/clk_out cp1_buffer1_0/clk_in cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs cp1_buffer1_2/charge_pump1_0/in7
+ VSUBS cp1_buffer1_2/vdd cp1_buffer1
Xcp1_buffer1_1 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_1/charge_pump1_0/vin
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_1/clk_out cp1_buffer1_1/clk_in cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs cp1_buffer1_2/charge_pump1_0/in7
+ VSUBS cp1_buffer1_2/vdd cp1_buffer1
Xcp1_buffer1_2 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/vin
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/clk_out cp1_buffer1_2/clk_in cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_2/charge_pump1_0/m1_12464_n576# cp1_buffer1_2/charge_pump1_0/in7 VSUBS
+ cp1_buffer1_2/vdd cp1_buffer1
Xcp1_buffer1_reverse_0 cp1_buffer1_1/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_1/clk_in
+ cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_2/vdd cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_0/clk_out
+ cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in7 VSUBS cp1_buffer1_reverse
Xcp1_buffer1_reverse_1 cp1_buffer1_2/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/clk_in
+ cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_2/vdd cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_1/clk_out
+ cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in7 VSUBS cp1_buffer1_reverse
C0 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in6 4.052151f
C1 cp1_buffer1_2/vdd cp1_buffer1_1/clk_out 2.547378f
C2 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in3 3.895406f
C3 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in2 3.972665f
C4 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in4 3.950372f
C5 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in7 3.640991f
C6 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in5 3.910277f
C7 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in1 4.003245f
C8 cp1_buffer1_2/vdd cp1_buffer1_0/clk_out 2.013929f
C9 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in8 3.700053f
C10 cp1_buffer1_2/vdd cp1_buffer1_1/clk_in 4.129703f
C11 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 VSUBS 22.596436f
C12 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C13 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C14 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C15 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C16 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C17 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C18 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C19 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C20 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C21 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C22 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C23 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C24 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_4341_n519# VSUBS 3.33176f
C25 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 VSUBS 22.21436f
C26 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_12659_300# VSUBS 2.683598f
C27 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C28 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C29 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C30 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C31 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C32 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C33 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C34 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C35 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C36 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C37 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C38 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C39 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C40 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C41 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C42 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C43 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C44 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C45 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C46 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C47 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C48 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C49 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C50 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C51 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C52 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C53 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C54 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C55 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C56 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C57 cp1_buffer1_2/charge_pump1_0/in8 VSUBS 11.267096f
C58 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C59 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk VSUBS 94.593094f
C60 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C61 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C62 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C63 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb VSUBS 0.101291p
C64 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C65 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C66 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2432_n962# VSUBS 8.68424f **FLOATING
C67 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2020_n482# VSUBS 2.56615f **FLOATING
C68 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_102# VSUBS 2.809951f
C69 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2402_572# VSUBS 2.172722f
C70 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_n986# VSUBS 2.381627f
C71 cp1_buffer1_2/clk_in VSUBS 7.486756f
C72 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_3246_118# VSUBS 6.834443f
C73 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 VSUBS 22.596436f
C74 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C75 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C76 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C77 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C78 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C79 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C80 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C81 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C82 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C83 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C84 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C85 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C86 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_4341_n519# VSUBS 3.33176f
C87 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 VSUBS 22.21436f
C88 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_12659_300# VSUBS 2.683598f
C89 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C90 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C91 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C92 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C93 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C94 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C95 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C96 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C97 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C98 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C99 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C100 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C101 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C102 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C103 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C104 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C105 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C106 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C107 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C108 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C109 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C110 cp1_buffer1_2/charge_pump1_0/in6 VSUBS 11.443146f
C111 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C112 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C113 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C114 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C115 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C116 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C117 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C118 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C119 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C120 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C121 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk VSUBS 94.698296f
C122 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C123 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C124 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C125 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb VSUBS 0.101284p
C126 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C127 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C128 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2432_n962# VSUBS 8.68424f **FLOATING
C129 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2020_n482# VSUBS 2.56615f **FLOATING
C130 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_102# VSUBS 2.809951f
C131 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2402_572# VSUBS 2.172722f
C132 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_n986# VSUBS 2.381627f
C133 cp1_buffer1_1/clk_in VSUBS 6.5659f
C134 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_3246_118# VSUBS 6.834443f
C135 cp1_buffer1_2/clk_out VSUBS 3.531028f
C136 cp1_buffer1_2/charge_pump1_0/input1 VSUBS 22.463037f
C137 cp1_buffer1_2/charge_pump1_0/input2 VSUBS 22.175997f
C138 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C139 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C140 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C141 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C142 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C143 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C144 cp1_buffer1_2/charge_pump1_0/in4 VSUBS 11.392217f
C145 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337917f
C146 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978384f
C147 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608259f
C148 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.339351f
C149 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.982591f
C150 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.609059f
C151 cp1_buffer1_2/charge_pump1_0/m1_4341_n519# VSUBS 3.771611f
C152 cp1_buffer1_2/charge_pump1_0/m1_12659_300# VSUBS 2.538747f
C153 cp1_buffer1_2/charge_pump1_0/m1_12464_n576# VSUBS 4.257501f
C154 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C155 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C156 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C157 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C158 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C159 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C160 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C161 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C162 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C163 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C164 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C165 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C166 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337823f
C167 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.9788f
C168 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608305f
C169 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337703f
C170 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978472f
C171 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608233f
C172 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C173 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C174 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C175 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C176 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C177 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C178 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.339689f
C179 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.984276f
C180 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.609388f
C181 cp1_buffer1_2/charge_pump1_0/in1 VSUBS 10.916974f
C182 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C183 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C184 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C185 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.3377f
C186 cp1_buffer1_2/charge_pump1_0/clkb VSUBS 89.72109f
C187 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.9784f
C188 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.608222f
C189 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C190 cp1_buffer1_2/charge_pump1_0/clk VSUBS 89.01907f
C191 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C192 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C193 cp1_buffer1_2/charge_pump1_0/clock_0/a_2432_n962# VSUBS 8.68424f **FLOATING
C194 cp1_buffer1_2/charge_pump1_0/clock_0/a_2020_n482# VSUBS 2.56615f **FLOATING
C195 cp1_buffer1_2/charge_pump1_0/clock_0/a_344_102# VSUBS 2.809951f
C196 cp1_buffer1_2/charge_pump1_0/clock_0/a_2402_572# VSUBS 2.172722f
C197 cp1_buffer1_2/charge_pump1_0/clock_0/a_344_n986# VSUBS 2.381627f
C198 cp1_buffer1_2/charge_pump1_0/clock_0/a_3246_118# VSUBS 6.834443f
C199 cp1_buffer1_2/charge_pump1_0/g2 VSUBS 2.344427f
C200 cp1_buffer1_2/charge_pump1_0/vin VSUBS 13.365224f
C201 cp1_buffer1_1/clk_out VSUBS 10.823749f
C202 cp1_buffer1_1/charge_pump1_0/input1 VSUBS 22.463037f
C203 cp1_buffer1_1/charge_pump1_0/input2 VSUBS 22.175129f
C204 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C205 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C206 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C207 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C208 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C209 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C210 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C211 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C212 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C213 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C214 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C215 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C216 cp1_buffer1_1/charge_pump1_0/m1_4341_n519# VSUBS 3.771611f
C217 cp1_buffer1_1/charge_pump1_0/m1_12659_300# VSUBS 2.538747f
C218 cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs VSUBS 14.537064f
C219 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C220 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C221 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C222 cp1_buffer1_2/charge_pump1_0/in7 VSUBS 10.908334f
C223 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C224 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C225 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C226 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C227 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C228 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C229 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C230 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C231 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C232 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C233 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C234 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C235 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C236 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C237 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C238 cp1_buffer1_2/charge_pump1_0/in2 VSUBS 11.33708f
C239 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C240 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C241 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C242 cp1_buffer1_2/charge_pump1_0/in3 VSUBS 11.200323f
C243 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C244 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C245 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C246 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C247 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C248 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C249 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C250 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C251 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C252 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C253 cp1_buffer1_1/charge_pump1_0/clkb VSUBS 89.843025f
C254 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C255 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C256 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C257 cp1_buffer1_1/charge_pump1_0/clk VSUBS 89.13844f
C258 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C259 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C260 cp1_buffer1_1/charge_pump1_0/clock_0/a_2432_n962# VSUBS 8.68424f **FLOATING
C261 cp1_buffer1_1/charge_pump1_0/clock_0/a_2020_n482# VSUBS 2.56615f **FLOATING
C262 cp1_buffer1_1/charge_pump1_0/clock_0/a_344_102# VSUBS 2.809951f
C263 cp1_buffer1_1/charge_pump1_0/clock_0/a_2402_572# VSUBS 2.172722f
C264 cp1_buffer1_1/charge_pump1_0/clock_0/a_344_n986# VSUBS 2.381627f
C265 cp1_buffer1_1/charge_pump1_0/clock_0/a_3246_118# VSUBS 6.834443f
C266 cp1_buffer1_1/charge_pump1_0/g2 VSUBS 2.344427f
C267 cp1_buffer1_1/charge_pump1_0/vin VSUBS 13.275853f
C268 cp1_buffer1_0/clk_in VSUBS 2.918218f
C269 cp1_buffer1_0/clk_out VSUBS 10.607181f
C270 cp1_buffer1_0/charge_pump1_0/input1 VSUBS 22.464737f
C271 cp1_buffer1_0/charge_pump1_0/input2 VSUBS 22.175129f
C272 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C273 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C274 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C275 cp1_buffer1_2/charge_pump1_0/in5 VSUBS 11.315837f
C276 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C277 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C278 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C279 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C280 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C281 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C282 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C283 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C284 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C285 cp1_buffer1_0/charge_pump1_0/m1_4341_n519# VSUBS 3.771611f
C286 cp1_buffer1_0/charge_pump1_0/m1_12659_300# VSUBS 2.538747f
C287 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs VSUBS 14.665705f
C288 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.340567f
C289 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.986715f
C290 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.609937f
C291 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.338885f
C292 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.980948f
C293 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608766f
C294 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.33837f
C295 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.979241f
C296 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608452f
C297 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C298 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C299 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C300 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C301 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C302 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C303 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C304 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C305 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C306 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C307 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C308 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C309 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337698f
C310 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978388f
C311 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C312 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C313 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C314 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C315 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.338463f
C316 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.979317f
C317 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608512f
C318 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C319 cp1_buffer1_0/charge_pump1_0/clkb VSUBS 89.82986f
C320 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C321 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
C322 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337703f
C323 cp1_buffer1_0/charge_pump1_0/clk VSUBS 88.92364f
C324 cp1_buffer1_2/vdd VSUBS 2.861079p
C325 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978397f
C326 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.608227f
C327 cp1_buffer1_0/charge_pump1_0/clock_0/a_2432_n962# VSUBS 8.68424f **FLOATING
C328 cp1_buffer1_0/charge_pump1_0/clock_0/a_2020_n482# VSUBS 2.56615f **FLOATING
C329 cp1_buffer1_0/charge_pump1_0/clock_0/a_344_102# VSUBS 2.809951f
C330 cp1_buffer1_0/charge_pump1_0/clock_0/a_2402_572# VSUBS 2.172722f
C331 cp1_buffer1_0/charge_pump1_0/clock_0/a_344_n986# VSUBS 2.381627f
C332 cp1_buffer1_0/charge_pump1_0/clock_0/a_3246_118# VSUBS 6.834443f
C333 cp1_buffer1_0/charge_pump1_0/g2 VSUBS 2.344427f
C334 cp1_buffer1_0/charge_pump1_0/vin VSUBS 10.37242f
.ends

.subckt sky130_fd_pr__nfet_01v8_D4CMYK a_15_n130# a_63_n42# a_n177_n130# a_255_n42#
+ a_n129_n42# a_111_64# a_n321_n42# a_159_n42# a_n81_64# a_n273_64# a_351_n42# a_207_n130#
+ a_303_64# a_n33_n42# a_n369_n130# a_n225_n42# a_n413_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_n130# a_n413_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt capacitor_5 cp_clk i1 vd2 vd1 vd4 vd3 clk GND VDD
Xbuffer_digital_1 i1 buffer_digital_1/in VDD GND buffer_digital
Xsky130_fd_pr__nfet_01v8_D4CMYK_0 vd2 GND vd2 GND GND vd2 GND GND vd2 vd2 GND vd2
+ vd2 GND vd2 GND GND GND sky130_fd_pr__nfet_01v8_D4CMYK
Xsky130_fd_pr__pfet_01v8_4ZKXAA_1 vd3 vd3 GND vd3 vd3 GND vd3 GND vd3 GND GND vd3
+ GND vd3 vd3 GND GND vd3 vd3 GND vd3 GND GND sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__pfet_01v8_4ZKXAA_2 vd4 vd4 GND vd4 vd4 GND vd4 GND vd4 GND GND vd4
+ GND vd4 vd4 GND GND vd4 vd4 GND vd4 GND GND sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__pfet_01v8_4ZKXAA_3 vd3 vd3 GND vd3 vd3 GND vd3 GND vd3 GND GND vd3
+ GND vd3 vd3 GND GND vd3 vd3 GND vd3 GND GND sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__nfet_01v8_NJGC45_0 GND vd1 GND vd1 vd1 GND GND vd1 vd1 GND vd1 GND
+ GND GND GND GND vd1 GND vd1 vd1 vd1 GND sky130_fd_pr__nfet_01v8_NJGC45
Xbuffer_and_gate_0 buffer_digital_1/in clk buffer_and_gate_0/out GND VDD buffer_and_gate
X0 buffer_and_gate_0/out cp_clk sky130_fd_pr__cap_mim_m3_1 l=4.97 w=5
C0 buffer_digital_1/in i1 2.935591f
C1 buffer_and_gate_0/and_gate_0/a_n78_396# GND 2.360761f
C2 clk GND 8.635434f
C3 VDD GND 20.988493f
C4 buffer_and_gate_0/buffer_0/a_1436_1552# GND 10.196393f
C5 vd1 GND 3.43263f
C6 vd3 GND 7.097779f
C7 vd4 GND 2.864619f
C8 vd2 GND 3.083021f
C9 buffer_digital_1/in GND 2.672912f
.ends

.subckt capacitors_5 capacitor_5_7/i1 capacitor_5_1/i1 capacitor_5_6/i1 capacitor_5_0/i1
+ capacitor_5_7/vd4 capacitor_5_3/i1 capacitor_5_7/vd2 capacitor_5_7/vd1 capacitor_5_7/cp_clk
+ capacitor_5_4/i1 capacitor_5_2/i1 capacitor_5_7/clk capacitor_5_7/vd3 capacitor_5_5/i1
+ VSUBS capacitor_5_7/VDD
Xcapacitor_5_5 capacitor_5_7/cp_clk capacitor_5_5/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_6 capacitor_5_7/cp_clk capacitor_5_6/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_7 capacitor_5_7/cp_clk capacitor_5_7/i1 capacitor_5_7/vd2 capacitor_5_7/vd1
+ capacitor_5_7/vd4 capacitor_5_7/vd3 capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_0 capacitor_5_7/cp_clk capacitor_5_0/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_1 capacitor_5_7/cp_clk capacitor_5_1/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_2 capacitor_5_7/cp_clk capacitor_5_2/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_3 capacitor_5_7/cp_clk capacitor_5_3/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_4 capacitor_5_7/cp_clk capacitor_5_4/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
C0 capacitor_5_7/VDD capacitor_5_7/cp_clk 11.685535f
C1 capacitor_5_7/VDD capacitor_5_7/clk 13.029696f
C2 capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.37575f
C3 capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.144792f
C4 capacitor_5_4/buffer_digital_1/in VSUBS 2.635156f
C5 capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.371064f
C6 capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.149221f
C7 capacitor_5_3/buffer_digital_1/in VSUBS 2.636791f
C8 capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.375672f
C9 capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.145726f
C10 capacitor_5_2/buffer_digital_1/in VSUBS 2.635774f
C11 capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.375235f
C12 capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.147629f
C13 capacitor_5_1/buffer_digital_1/in VSUBS 2.636666f
C14 capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C15 capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C16 capacitor_5_0/buffer_digital_1/in VSUBS 2.58165f
C17 capacitor_5_7/cp_clk VSUBS 20.068026f
C18 capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.376815f
C19 capacitor_5_7/clk VSUBS 71.174866f
C20 capacitor_5_7/VDD VSUBS 0.260321p
C21 capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.147582f
C22 capacitor_5_7/vd1 VSUBS 2.321869f
C23 capacitor_5_7/vd3 VSUBS 3.828029f
C24 capacitor_5_7/vd2 VSUBS 2.223177f
C25 capacitor_5_7/buffer_digital_1/in VSUBS 2.636351f
C26 capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.376023f
C27 capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.14572f
C28 capacitor_5_6/buffer_digital_1/in VSUBS 2.635363f
C29 capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.376738f
C30 capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.148531f
C31 capacitor_5_5/buffer_digital_1/in VSUBS 2.636503f
.ends

.subckt nmos_diode2 a_350_n764# a_970_n762# a_410_n892# dw_118_n1078# VSUBS
X0 a_410_n892# a_410_n892# a_350_n764# dw_118_n1078# sky130_fd_pr__nfet_01v8 ad=0.8729 pd=6.6 as=0.9029 ps=6.62 w=3.01 l=1
X1 a_350_n764# a_970_n762# a_970_n762# dw_118_n1078# sky130_fd_pr__nfet_01v8 ad=0.9929 pd=6.68 as=0.8729 ps=6.6 w=3.01 l=1
C0 dw_118_n1078# VSUBS 8.163819f
.ends

.subckt charge_pump in1 in3 in5 input1 input2 out clk clkb clk_in g1 g2 vin a_18057_18271#
+ in6 in8 in4 in7 in2 vs clock_0/gnd clock_0/vdd
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 g1 clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 g2 clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xcapacitors_5_1 in8 in2 in7 in1 clock_0/vdd in4 clock_0/vdd clock_0/vdd input2 in5
+ in3 clkb clock_0/vdd in6 clock_0/gnd clock_0/vdd capacitors_5
Xcapacitors_5_0 in8 in2 in7 in1 clock_0/vdd in4 clock_0/vdd clock_0/vdd input1 in5
+ in3 clk clock_0/vdd in6 clock_0/gnd clock_0/vdd capacitors_5
Xnmos_dnw3_0 vin input1 input2 g1 g2 vs clock_0/gnd nmos_dnw3
Xclock_0 clk_in clock_0/vdd clock_0/gnd clk clkb clock
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xnmos_diode2_0 out input2 input1 vs nmos_diode2_0/VSUBS nmos_diode2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 input2 clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 input1 clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 vs clkb 2.334149f
C1 clock_0/vdd vs 11.967723f
C2 vs input2 4.024266f
C3 clock_0/vdd clkb 17.402271f
C4 clk vs 2.642354f
C5 out vs 14.162663f
C6 clock_0/vdd clk 26.498405f
C7 out clock_0/vdd 2.310455f
C8 input1 vs 3.387235f
C9 vs vin 8.809598f
C10 input1 input2 8.763355f
C11 clock_0/vdd vin 5.355844f
C12 vs nmos_diode2_0/VSUBS 20.067162f
C13 out nmos_diode2_0/VSUBS 3.142924f
C14 clock_0/a_2432_n962# nmos_diode2_0/VSUBS 8.684403f **FLOATING
C15 clock_0/a_2020_n482# nmos_diode2_0/VSUBS 2.571413f **FLOATING
C16 clock_0/a_344_102# nmos_diode2_0/VSUBS 2.810446f
C17 clock_0/a_2402_572# nmos_diode2_0/VSUBS 2.172722f
C18 clock_0/a_344_n986# nmos_diode2_0/VSUBS 2.381627f
C19 clock_0/a_3246_118# nmos_diode2_0/VSUBS 6.834443f
C20 g2 nmos_diode2_0/VSUBS 2.43748f
C21 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C22 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978447f
C23 capacitors_5_0/capacitor_5_4/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581751f
C24 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C25 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C26 capacitors_5_0/capacitor_5_3/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581653f
C27 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C28 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C29 capacitors_5_0/capacitor_5_2/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C30 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C31 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C32 capacitors_5_0/capacitor_5_1/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C33 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C34 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978566f
C35 capacitors_5_0/capacitor_5_0/buffer_digital_1/in nmos_diode2_0/VSUBS 2.583461f
C36 input1 nmos_diode2_0/VSUBS 16.681173f
C37 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C38 clk nmos_diode2_0/VSUBS 84.957054f
C39 clock_0/vdd nmos_diode2_0/VSUBS 0.459957p
C40 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978453f
C41 capacitors_5_0/capacitor_5_7/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581764f
C42 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C43 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978465f
C44 capacitors_5_0/capacitor_5_6/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581762f
C45 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C46 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978452f
C47 capacitors_5_0/capacitor_5_5/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581756f
C48 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C49 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C50 capacitors_5_1/capacitor_5_4/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C51 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C52 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.97846f
C53 capacitors_5_1/capacitor_5_3/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581745f
C54 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C55 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978502f
C56 capacitors_5_1/capacitor_5_2/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581764f
C57 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C58 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978491f
C59 capacitors_5_1/capacitor_5_1/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58176f
C60 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C61 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978744f
C62 capacitors_5_1/capacitor_5_0/buffer_digital_1/in nmos_diode2_0/VSUBS 2.583578f
C63 input2 nmos_diode2_0/VSUBS 16.89145f
C64 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C65 clkb nmos_diode2_0/VSUBS 87.08427f
C66 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C67 capacitors_5_1/capacitor_5_7/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581653f
C68 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C69 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C70 capacitors_5_1/capacitor_5_6/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C71 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C72 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C73 capacitors_5_1/capacitor_5_5/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C74 g1 nmos_diode2_0/VSUBS 2.639545f
.ends

.subckt cp2_buffer1 charge_pump_0/a_18057_18271# charge_pump_0/in4 buffer_digital_0/in
+ charge_pump_0/in5 charge_pump_0/vin charge_pump_0/out charge_pump_0/in6 charge_pump_0/in7
+ charge_pump_0/vs charge_pump_0/in8 charge_pump_0/in1 charge_pump_0/in3 charge_pump_0/in2
+ buffer_digital_1/i VSUBS buffer_digital_1/VDD
Xpmos_decap_10_10 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_11 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_12 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_13 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xcharge_pump_0 charge_pump_0/in1 charge_pump_0/in3 charge_pump_0/in5 charge_pump_0/input1
+ charge_pump_0/input2 charge_pump_0/out charge_pump_0/clk charge_pump_0/clkb buffer_digital_0/in
+ charge_pump_0/g1 charge_pump_0/g2 charge_pump_0/vin charge_pump_0/a_18057_18271#
+ charge_pump_0/in6 charge_pump_0/in8 charge_pump_0/in4 charge_pump_0/in7 charge_pump_0/in2
+ charge_pump_0/vs VSUBS buffer_digital_1/VDD charge_pump
Xbuffer_digital_0 buffer_digital_0/i buffer_digital_0/in buffer_digital_1/VDD VSUBS
+ buffer_digital
Xbuffer_digital_1 buffer_digital_1/i buffer_digital_0/i buffer_digital_1/VDD VSUBS
+ buffer_digital
Xnmos_decap_10_0 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_1 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_2 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_3 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_4 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_5 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_0 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_1 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_2 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_3 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_4 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_5 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_6 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_7 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_9 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_8 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
C0 buffer_digital_0/in buffer_digital_1/VDD 4.800197f
C1 buffer_digital_1/VDD buffer_digital_1/i 3.73526f
C2 buffer_digital_1/i charge_pump_0/nmos_diode2_0/VSUBS 8.29284f
C3 charge_pump_0/vs charge_pump_0/nmos_diode2_0/VSUBS 18.969007f
C4 charge_pump_0/clock_0/a_2432_n962# charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C5 charge_pump_0/clock_0/a_2020_n482# charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C6 charge_pump_0/clock_0/a_344_102# charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C7 charge_pump_0/clock_0/a_2402_572# charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C8 charge_pump_0/clock_0/a_344_n986# charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C9 buffer_digital_0/in charge_pump_0/nmos_diode2_0/VSUBS 12.889783f
C10 charge_pump_0/clock_0/a_3246_118# charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C11 charge_pump_0/g2 charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C12 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C13 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C14 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C15 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C16 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C17 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C18 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C19 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C20 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C21 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C22 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C23 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C24 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C25 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C26 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C27 charge_pump_0/input1 charge_pump_0/nmos_diode2_0/VSUBS 15.031953f
C28 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C29 charge_pump_0/clk charge_pump_0/nmos_diode2_0/VSUBS 82.80111f
C30 buffer_digital_1/VDD charge_pump_0/nmos_diode2_0/VSUBS 0.525238p
C31 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C32 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C33 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C34 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C35 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C36 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C37 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C38 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C39 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C40 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C41 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C42 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C43 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C44 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C45 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C46 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C47 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C48 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C49 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C50 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C51 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C52 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C53 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C54 charge_pump_0/input2 charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C55 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C56 charge_pump_0/clkb charge_pump_0/nmos_diode2_0/VSUBS 83.927444f
C57 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C58 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C59 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C60 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C61 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C62 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C63 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C64 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C65 charge_pump_0/g1 charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
.ends

.subckt charge_pump_reverse m1_11946_n452# nmos_dnw3_0/vin capacitors_5_1/capacitor_5_2/i1
+ capacitors_5_1/capacitor_5_3/i1 a_18057_18271# capacitors_5_1/capacitor_5_4/i1 capacitors_5_1/capacitor_5_5/i1
+ clock_0/clk_in clock_0/vdd capacitors_5_1/capacitor_5_0/i1 capacitors_5_1/capacitor_5_7/i1
+ clock_0/gnd capacitors_5_1/capacitor_5_6/i1 capacitors_5_1/capacitor_5_1/i1 nmos_dnw3_0/vs
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xcapacitors_5_1 capacitors_5_1/capacitor_5_7/i1 capacitors_5_1/capacitor_5_1/i1 capacitors_5_1/capacitor_5_6/i1
+ capacitors_5_1/capacitor_5_0/i1 clock_0/vdd capacitors_5_1/capacitor_5_3/i1 clock_0/vdd
+ clock_0/vdd nmos_dnw3_0/out2 capacitors_5_1/capacitor_5_4/i1 capacitors_5_1/capacitor_5_2/i1
+ clock_0/clk clock_0/vdd capacitors_5_1/capacitor_5_5/i1 clock_0/gnd clock_0/vdd
+ capacitors_5
Xcapacitors_5_0 capacitors_5_1/capacitor_5_7/i1 capacitors_5_1/capacitor_5_1/i1 capacitors_5_1/capacitor_5_6/i1
+ capacitors_5_1/capacitor_5_0/i1 clock_0/vdd capacitors_5_1/capacitor_5_3/i1 clock_0/vdd
+ clock_0/vdd nmos_dnw3_0/out1 capacitors_5_1/capacitor_5_4/i1 capacitors_5_1/capacitor_5_2/i1
+ clock_0/clkb clock_0/vdd capacitors_5_1/capacitor_5_5/i1 clock_0/gnd clock_0/vdd
+ capacitors_5
Xnmos_dnw3_0 nmos_dnw3_0/vin nmos_dnw3_0/out1 nmos_dnw3_0/out2 nmos_dnw3_0/clk nmos_dnw3_0/clkb
+ nmos_dnw3_0/vs clock_0/gnd nmos_dnw3
Xclock_0 clock_0/clk_in clock_0/vdd clock_0/gnd clock_0/clk clock_0/clkb clock
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xnmos_diode2_0 m1_11946_n452# nmos_dnw3_0/out2 nmos_dnw3_0/out1 nmos_dnw3_0/vs clock_0/gnd
+ nmos_diode2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 nmos_dnw3_0/out2 clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 nmos_dnw3_0/out1 clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 clock_0/vdd nmos_dnw3_0/vs 2.471132f
C1 m1_11946_n452# nmos_dnw3_0/vs 13.479089f
C2 clock_0/vdd m1_11946_n452# 2.540002f
C3 nmos_dnw3_0/out2 nmos_dnw3_0/out1 8.763353f
C4 nmos_dnw3_0/out1 nmos_dnw3_0/vs 3.314235f
C5 clock_0/clkb clock_0/vdd 24.445723f
C6 clock_0/vdd clock_0/clk 20.032824f
C7 nmos_dnw3_0/vin clock_0/vdd 8.882092f
C8 nmos_dnw3_0/out2 nmos_dnw3_0/vs 5.257541f
C9 nmos_dnw3_0/vs clock_0/gnd 19.463373f
C10 m1_11946_n452# clock_0/gnd 2.969539f
C11 clock_0/a_2432_n962# clock_0/gnd 8.689615f **FLOATING
C12 clock_0/a_2020_n482# clock_0/gnd 2.568188f **FLOATING
C13 clock_0/a_344_102# clock_0/gnd 2.809951f
C14 clock_0/a_2402_572# clock_0/gnd 2.172722f
C15 clock_0/a_344_n986# clock_0/gnd 2.381627f
C16 clock_0/a_3246_118# clock_0/gnd 6.834443f
C17 nmos_dnw3_0/vin clock_0/gnd 2.49859f
C18 nmos_dnw3_0/clkb clock_0/gnd 2.242713f
C19 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C20 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978447f
C21 capacitors_5_0/capacitor_5_4/buffer_digital_1/in clock_0/gnd 2.581751f
C22 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C23 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C24 capacitors_5_0/capacitor_5_3/buffer_digital_1/in clock_0/gnd 2.581652f
C25 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C26 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C27 capacitors_5_0/capacitor_5_2/buffer_digital_1/in clock_0/gnd 2.581652f
C28 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C29 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C30 capacitors_5_0/capacitor_5_1/buffer_digital_1/in clock_0/gnd 2.581652f
C31 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C32 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978566f
C33 capacitors_5_0/capacitor_5_0/buffer_digital_1/in clock_0/gnd 2.583461f
C34 nmos_dnw3_0/out1 clock_0/gnd 16.704819f
C35 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C36 clock_0/clkb clock_0/gnd 92.38439f
C37 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978453f
C38 capacitors_5_0/capacitor_5_7/buffer_digital_1/in clock_0/gnd 2.581764f
C39 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C40 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978465f
C41 capacitors_5_0/capacitor_5_6/buffer_digital_1/in clock_0/gnd 2.581762f
C42 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C43 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978452f
C44 capacitors_5_0/capacitor_5_5/buffer_digital_1/in clock_0/gnd 2.581756f
C45 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C46 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C47 capacitors_5_1/capacitor_5_4/buffer_digital_1/in clock_0/gnd 2.581652f
C48 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C49 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.97846f
C50 capacitors_5_1/capacitor_5_3/buffer_digital_1/in clock_0/gnd 2.581745f
C51 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C52 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978502f
C53 capacitors_5_1/capacitor_5_2/buffer_digital_1/in clock_0/gnd 2.581763f
C54 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C55 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978491f
C56 capacitors_5_1/capacitor_5_1/buffer_digital_1/in clock_0/gnd 2.58176f
C57 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C58 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978744f
C59 capacitors_5_1/capacitor_5_0/buffer_digital_1/in clock_0/gnd 2.583578f
C60 nmos_dnw3_0/out2 clock_0/gnd 16.02703f
C61 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C62 clock_0/clk clock_0/gnd 86.04303f
C63 clock_0/vdd clock_0/gnd 0.45817p
C64 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C65 capacitors_5_1/capacitor_5_7/buffer_digital_1/in clock_0/gnd 2.581653f
C66 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C67 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C68 capacitors_5_1/capacitor_5_6/buffer_digital_1/in clock_0/gnd 2.581652f
C69 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C70 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C71 capacitors_5_1/capacitor_5_5/buffer_digital_1/in clock_0/gnd 2.581652f
C72 nmos_dnw3_0/clk clock_0/gnd 2.52759f
.ends

.subckt cp2_buffer2 buffer_digital_3/in charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/i1
+ charge_pump_reverse_0/nmos_dnw3_0/vin charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/i1
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/i1 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/i1
+ buffer_digital_3/VDD charge_pump_reverse_0/nmos_dnw3_0/vs charge_pump_reverse_0/m1_11946_n452#
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/i1 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/i1
+ buffer_digital_2/i charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/i1 VSUBS charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/i1
Xpmos_decap_10_10 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_11 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_12 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_13 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_14 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_15 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xbuffer_digital_2 buffer_digital_2/i buffer_digital_3/i buffer_digital_3/VDD VSUBS
+ buffer_digital
Xbuffer_digital_3 buffer_digital_3/i buffer_digital_3/in buffer_digital_3/VDD VSUBS
+ buffer_digital
Xnmos_decap_10_0 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_1 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xcharge_pump_reverse_0 charge_pump_reverse_0/m1_11946_n452# charge_pump_reverse_0/nmos_dnw3_0/vin
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/i1 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/i1
+ VSUBS charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/i1 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/i1
+ buffer_digital_3/in buffer_digital_3/VDD charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/i1
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/i1 VSUBS charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/i1
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/i1 charge_pump_reverse_0/nmos_dnw3_0/vs
+ charge_pump_reverse
Xnmos_decap_10_2 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_3 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_4 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_5 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_6 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_7 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_8 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_9 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_0 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_1 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_2 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_3 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_4 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_5 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_6 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_7 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_9 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_8 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
C0 buffer_digital_3/VDD buffer_digital_2/i 3.650215f
C1 buffer_digital_3/VDD buffer_digital_3/in 5.148005f
C2 charge_pump_reverse_0/clock_0/clkb buffer_digital_3/VDD 3.552189f
C3 charge_pump_reverse_0/nmos_dnw3_0/vs VSUBS 18.79532f
C4 charge_pump_reverse_0/clock_0/a_2432_n962# VSUBS 8.68424f **FLOATING
C5 charge_pump_reverse_0/clock_0/a_2020_n482# VSUBS 2.56615f **FLOATING
C6 charge_pump_reverse_0/clock_0/a_344_102# VSUBS 2.809951f
C7 charge_pump_reverse_0/clock_0/a_2402_572# VSUBS 2.172722f
C8 charge_pump_reverse_0/clock_0/a_344_n986# VSUBS 2.381627f
C9 buffer_digital_3/in VSUBS 11.44915f
C10 charge_pump_reverse_0/clock_0/a_3246_118# VSUBS 6.834443f
C11 charge_pump_reverse_0/nmos_dnw3_0/vin VSUBS 2.458278f
C12 charge_pump_reverse_0/nmos_dnw3_0/clkb VSUBS 2.234749f
C13 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C14 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C15 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in VSUBS 2.581652f
C16 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C17 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C18 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in VSUBS 2.581652f
C19 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C20 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C21 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in VSUBS 2.581652f
C22 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C23 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C24 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in VSUBS 2.581652f
C25 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C26 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C27 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in VSUBS 2.581652f
C28 charge_pump_reverse_0/nmos_dnw3_0/out1 VSUBS 15.064581f
C29 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C30 charge_pump_reverse_0/clock_0/clkb VSUBS 90.50171f
C31 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C32 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in VSUBS 2.581652f
C33 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C34 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C35 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in VSUBS 2.581652f
C36 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C37 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C38 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in VSUBS 2.581652f
C39 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C40 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C41 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in VSUBS 2.581652f
C42 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C43 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C44 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in VSUBS 2.581652f
C45 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C46 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C47 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in VSUBS 2.581652f
C48 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C49 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C50 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in VSUBS 2.581652f
C51 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C52 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C53 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in VSUBS 2.581652f
C54 charge_pump_reverse_0/nmos_dnw3_0/out2 VSUBS 14.843945f
C55 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C56 charge_pump_reverse_0/clock_0/clk VSUBS 84.616936f
C57 buffer_digital_3/VDD VSUBS 0.546588p
C58 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C59 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in VSUBS 2.581652f
C60 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C61 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C62 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in VSUBS 2.581652f
C63 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C64 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C65 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in VSUBS 2.581652f
C66 charge_pump_reverse_0/nmos_dnw3_0/clk VSUBS 2.425359f
C67 buffer_digital_2/i VSUBS 10.683858f
.ends

.subckt cp2_buffer_5stage cp2_buffer1_0/charge_pump_0/vin cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer1_1/charge_pump_0/out cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer1_2/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_0/charge_pump_0/out
+ cp2_buffer1_2/charge_pump_0/in3 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/vs
+ cp2_buffer1_1/charge_pump_0/vs cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/vs
+ cp2_buffer1_2/charge_pump_0/in4 cp2_buffer1_2/charge_pump_0/out cp2_buffer1_2/buffer_digital_0/in
+ cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/in7 cp2_buffer1_0/charge_pump_0/vs
+ cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_0/buffer_digital_1/i
+ cp2_buffer1_2/charge_pump_0/a_18057_18271# VSUBS
Xcp2_buffer1_0 cp2_buffer1_0/charge_pump_0/a_18057_18271# cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer2_0/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_0/charge_pump_0/vin
+ cp2_buffer1_0/charge_pump_0/out cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in7
+ cp2_buffer1_0/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_0/buffer_digital_1/i
+ VSUBS cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1
Xcp2_buffer1_1 cp2_buffer1_1/charge_pump_0/a_18057_18271# cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer2_1/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer1_1/charge_pump_0/out cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in7
+ cp2_buffer1_1/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_1/buffer_digital_1/i
+ VSUBS cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1
Xcp2_buffer1_2 cp2_buffer1_2/charge_pump_0/a_18057_18271# cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer1_2/buffer_digital_0/in cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/vin
+ cp2_buffer1_2/charge_pump_0/out cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in7
+ cp2_buffer1_2/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_2/buffer_digital_1/i
+ VSUBS cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1
Xcp2_buffer2_0 cp2_buffer1_1/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/in7 cp2_buffer1_0/charge_pump_0/out
+ cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/vs
+ cp2_buffer1_1/charge_pump_0/vin cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer2_0/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/in8 VSUBS cp2_buffer1_2/charge_pump_0/in2
+ cp2_buffer2
Xcp2_buffer2_1 cp2_buffer1_2/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/in7 cp2_buffer1_1/charge_pump_0/out
+ cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/vs
+ cp2_buffer1_2/charge_pump_0/vin cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer2_1/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/in8 VSUBS cp2_buffer1_2/charge_pump_0/in2
+ cp2_buffer2
C0 cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/in2 4.401648f
C1 cp2_buffer1_2/charge_pump_0/in4 cp2_buffer2_1/buffer_digital_3/VDD 4.388158f
C2 cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/in8 4.645438f
C3 cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/in5 4.394f
C4 cp2_buffer1_2/charge_pump_0/in1 cp2_buffer2_1/buffer_digital_3/VDD 4.323198f
C5 cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/in6 4.452658f
C6 cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/in3 4.418769f
C7 cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/in7 4.44695f
C8 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 18.79948f
C9 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C10 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C11 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C12 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C13 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C14 cp2_buffer1_2/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.964601f
C15 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C16 cp2_buffer1_1/charge_pump_0/out cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.876493f
C17 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.234749f
C18 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C19 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C20 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C21 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C22 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C23 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C24 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C25 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C26 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C27 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C28 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C29 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C30 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C31 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C32 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C33 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.064581f
C34 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C35 cp2_buffer2_1/charge_pump_reverse_0/clock_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.96087f
C36 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C37 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C38 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C39 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C40 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C41 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C42 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C43 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C44 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C45 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C46 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C47 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C48 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C49 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C50 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C51 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C52 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C53 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C54 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C55 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C56 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C57 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C58 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C59 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.843945f
C60 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C61 cp2_buffer2_1/charge_pump_reverse_0/clock_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.546394f
C62 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C63 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C64 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C65 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C66 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C67 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C68 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C69 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C70 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.425359f
C71 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 18.799305f
C72 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C73 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C74 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C75 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C76 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C77 cp2_buffer1_1/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.7906f
C78 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C79 cp2_buffer1_0/charge_pump_0/out cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 4.363251f
C80 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.234749f
C81 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C82 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C83 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C84 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C85 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C86 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C87 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C88 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C89 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C90 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C91 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C92 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C93 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C94 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C95 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C96 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.064581f
C97 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C98 cp2_buffer2_0/charge_pump_reverse_0/clock_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.90249f
C99 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C100 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C101 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C102 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C103 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C104 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C105 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C106 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C107 cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.731117f
C108 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C109 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C110 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C111 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C112 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C113 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C114 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C115 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C116 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C117 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C118 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C119 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C120 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C121 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C122 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C123 cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.184977f
C124 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.843945f
C125 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C126 cp2_buffer2_0/charge_pump_reverse_0/clock_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.56565f
C127 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C128 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C129 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C130 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C131 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C132 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C133 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C134 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C135 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.425359f
C136 cp2_buffer1_2/charge_pump_0/vin cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.491769f
C137 cp2_buffer1_2/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 18.960741f
C138 cp2_buffer1_2/charge_pump_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C139 cp2_buffer1_2/charge_pump_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C140 cp2_buffer1_2/charge_pump_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C141 cp2_buffer1_2/charge_pump_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C142 cp2_buffer1_2/charge_pump_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C143 cp2_buffer1_2/buffer_digital_0/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 4.599239f
C144 cp2_buffer1_2/charge_pump_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C145 cp2_buffer1_2/charge_pump_0/g2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C146 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C147 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C148 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C149 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C150 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C151 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C152 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C153 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C154 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C155 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C156 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C157 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C158 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C159 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C160 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C161 cp2_buffer1_2/charge_pump_0/input1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.031953f
C162 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C163 cp2_buffer1_2/charge_pump_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.45232f
C164 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C165 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C166 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C167 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C168 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C169 cp2_buffer1_2/charge_pump_0/in7 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.785422f
C170 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C171 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C172 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C173 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C174 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C175 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C176 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C177 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C178 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C179 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C180 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C181 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C182 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C183 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C184 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C185 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C186 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C187 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C188 cp2_buffer1_2/charge_pump_0/input2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C189 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C190 cp2_buffer1_2/charge_pump_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.803345f
C191 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C192 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C193 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C194 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C195 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C196 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C197 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C198 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C199 cp2_buffer1_2/charge_pump_0/g1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
C200 cp2_buffer1_1/charge_pump_0/vin cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.621271f
C201 cp2_buffer1_1/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 18.970835f
C202 cp2_buffer1_1/charge_pump_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C203 cp2_buffer1_1/charge_pump_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C204 cp2_buffer1_1/charge_pump_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C205 cp2_buffer1_1/charge_pump_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C206 cp2_buffer1_1/charge_pump_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C207 cp2_buffer2_1/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.156822f
C208 cp2_buffer1_1/charge_pump_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C209 cp2_buffer1_1/charge_pump_0/g2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C210 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C211 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C212 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C213 cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.690011f
C214 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C215 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C216 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C217 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C218 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C219 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C220 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C221 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C222 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C223 cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.795872f
C224 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C225 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C226 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C227 cp2_buffer1_1/charge_pump_0/input1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.031953f
C228 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C229 cp2_buffer1_1/charge_pump_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.48422f
C230 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C231 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C232 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C233 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C234 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C235 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C236 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C237 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C238 cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.70006f
C239 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C240 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C241 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C242 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C243 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C244 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C245 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C246 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C247 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C248 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C249 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C250 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C251 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C252 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C253 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C254 cp2_buffer1_1/charge_pump_0/input2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C255 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C256 cp2_buffer1_1/charge_pump_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.94922f
C257 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C258 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C259 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C260 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C261 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C262 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C263 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C264 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C265 cp2_buffer1_1/charge_pump_0/g1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
C266 cp2_buffer1_0/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 4.024008f
C267 cp2_buffer1_0/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 18.96282f
C268 cp2_buffer1_0/charge_pump_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C269 cp2_buffer1_0/charge_pump_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C270 cp2_buffer1_0/charge_pump_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C271 cp2_buffer1_0/charge_pump_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C272 cp2_buffer1_0/charge_pump_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C273 cp2_buffer2_0/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.215527f
C274 cp2_buffer1_0/charge_pump_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C275 cp2_buffer1_0/charge_pump_0/g2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C276 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337914f
C277 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.977524f
C278 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58151f
C279 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337862f
C280 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.979101f
C281 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581781f
C282 cp2_buffer1_2/charge_pump_0/in4 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.693232f
C283 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.338461f
C284 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.981709f
C285 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.582303f
C286 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337865f
C287 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.97974f
C288 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581686f
C289 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337563f
C290 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978114f
C291 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581487f
C292 cp2_buffer1_2/charge_pump_0/in1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.087496f
C293 cp2_buffer1_0/charge_pump_0/input1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.034381f
C294 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.340502f
C295 cp2_buffer1_0/charge_pump_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.13737f
C296 cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.562668p
C297 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.985868f
C298 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.583144f
C299 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337697f
C300 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978412f
C301 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C302 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.339153f
C303 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.981775f
C304 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.582313f
C305 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C306 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C307 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C308 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C309 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C310 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C311 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C312 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C313 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C314 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C315 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C316 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C317 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C318 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C319 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C320 cp2_buffer1_0/charge_pump_0/input2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C321 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C322 cp2_buffer1_0/charge_pump_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.94053f
C323 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C324 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C325 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C326 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C327 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C328 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C329 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C330 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C331 cp2_buffer1_0/charge_pump_0/g1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
.ends

.subckt reconfigurable_CP1
Xcp1_buffer_5stage_0 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in8
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in7 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in6
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in5
+ cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vin cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer_5stage_0/cp1_buffer1_0/clk_in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in4
+ cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/vin cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/vin
+ cp1_buffer_5stage_0/cp1_buffer1_2/vdd VSUBS cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in3
+ cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vs cp1_buffer_5stage
Xcp2_buffer_5stage_0 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in8 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vs
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in7 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vs
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in6 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vin
+ cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vs cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in5 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vin
+ cp2_buffer_5stage_0/cp2_buffer1_2/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in2 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vs
+ cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in3
+ cp2_buffer_5stage_0/cp2_buffer1_0/buffer_digital_1/i cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/a_18057_18271#
+ VSUBS cp2_buffer_5stage
Xcp2_buffer_5stage_1 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in8
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/vs
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in2 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vs
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in3 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vin
+ cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in4 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/out
+ cp2_buffer_5stage_0/cp2_buffer1_0/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in5
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in7 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vs
+ cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in6
+ cp1_buffer_5stage_0/cp1_buffer1_0/clk_in VSUBS VSUBS cp2_buffer_5stage
C0 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in6 3.297943f
C1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in7 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in3 2.23645f
C2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in5 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in4 10.4178f
C3 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in7 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in6 8.12519f
C4 cp1_buffer_5stage_0/cp1_buffer1_0/clk_in cp1_buffer_5stage_0/cp1_buffer1_2/vdd 9.963273f
C5 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in7 3.749474f
C6 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in5 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in6 9.032085f
C7 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in1 2.384012f
C8 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_0/cp2_buffer1_0/buffer_digital_1/i 8.525254f
C9 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in5 3.039896f
C10 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in3 8.1524f
C11 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in8 3.171637f
C12 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in4 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in3 9.04317f
C13 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in7 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in8 5.25029f
C14 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in2 2.844454f
C15 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in8 3.24343f
C16 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in4 2.62203f
C17 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in3 2.54084f
C18 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in7 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in2 2.68839f
C19 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in2 13.281401f
C20 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 23.166407f
C21 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C22 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C23 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C24 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C25 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C26 cp2_buffer_5stage_1/cp2_buffer1_2/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.412422f
C27 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C28 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.234749f
C29 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C30 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C31 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C32 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C33 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C34 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C35 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C36 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C37 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C38 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C39 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C40 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C41 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C42 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C43 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C44 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.064581f
C45 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C46 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.91548f
C47 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C48 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C49 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C50 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C51 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C52 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C53 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C54 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C55 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C56 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C57 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C58 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C59 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C60 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C61 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C62 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C63 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C64 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C65 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C66 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C67 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C68 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C69 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C70 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.843945f
C71 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C72 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.49679f
C73 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C74 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C75 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C76 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C77 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C78 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C79 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C80 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C81 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.425359f
C82 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 28.936113f
C83 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C84 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C85 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C86 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C87 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C88 cp2_buffer_5stage_1/cp2_buffer1_1/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.267972f
C89 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C90 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.234749f
C91 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C92 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C93 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C94 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C95 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C96 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C97 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C98 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C99 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C100 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C101 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C102 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C103 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C104 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C105 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C106 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.064581f
C107 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C108 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.91548f
C109 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C110 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C111 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C112 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C113 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C114 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C115 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C116 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C117 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in3 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 36.902527f
C118 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C119 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C120 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C121 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C122 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C123 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C124 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C125 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C126 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C127 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C128 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C129 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C130 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C131 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C132 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C133 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in8 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 56.946053f
C134 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.843945f
C135 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C136 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.49679f
C137 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C138 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C139 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C140 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C141 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C142 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C143 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C144 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C145 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.425359f
C146 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.284825f
C147 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 23.301306f
C148 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C149 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C150 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C151 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C152 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C153 cp2_buffer_5stage_0/cp2_buffer1_0/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 11.466456f
C154 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C155 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C156 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C157 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C158 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C159 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C160 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C161 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C162 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C163 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C164 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C165 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C166 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C167 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C168 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C169 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C170 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C171 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.031953f
C172 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C173 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.29479f
C174 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C175 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C176 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C177 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C178 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C179 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C180 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C181 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C182 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C183 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C184 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C185 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C186 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C187 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C188 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C189 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C190 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C191 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C192 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C193 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C194 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C195 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C196 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C197 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C198 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C199 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.85823f
C200 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C201 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C202 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C203 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C204 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C205 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C206 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C207 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C208 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
C209 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 24.129698f
C210 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C211 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C212 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C213 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C214 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C215 cp2_buffer_5stage_1/cp2_buffer2_1/buffer_digital_2/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.84415f
C216 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C217 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C218 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C219 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C220 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C221 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C222 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C223 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C224 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C225 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C226 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C227 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C228 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C229 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C230 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 35.499798f
C231 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C232 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C233 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C234 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.031953f
C235 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C236 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.29458f
C237 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C238 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C239 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C240 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C241 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C242 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C243 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C244 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C245 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in6 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 30.626343f
C246 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C247 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C248 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C249 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C250 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C251 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C252 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C253 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C254 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C255 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C256 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C257 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C258 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C259 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C260 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C261 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C262 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C263 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.97966f
C264 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C265 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C266 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C267 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C268 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C269 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C270 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C271 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C272 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
C273 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 50.312313f
C274 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C275 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C276 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C277 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C278 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C279 cp2_buffer_5stage_1/cp2_buffer2_0/buffer_digital_2/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.985027f
C280 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C281 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C282 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C283 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C284 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C285 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C286 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C287 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C288 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in4 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 35.164486f
C289 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C290 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C291 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C292 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C293 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C294 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C295 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C296 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C297 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C298 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.031953f
C299 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C300 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.243904f
C301 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C302 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C303 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C304 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C305 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C306 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C307 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C308 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C309 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C310 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C311 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C312 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C313 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C314 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C315 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C316 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C317 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C318 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C319 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C320 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C321 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C322 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C323 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C324 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C325 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C326 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.97966f
C327 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C328 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C329 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C330 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C331 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C332 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C333 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C334 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C335 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
C336 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 23.114765f
C337 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C338 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C339 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C340 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C341 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C342 cp2_buffer_5stage_0/cp2_buffer1_2/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.371514f
C343 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C344 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.234749f
C345 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C346 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C347 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C348 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C349 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C350 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C351 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C352 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C353 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C354 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C355 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C356 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C357 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C358 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C359 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C360 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.064581f
C361 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C362 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.91548f
C363 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C364 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C365 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C366 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C367 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C368 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C369 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C370 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C371 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C372 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C373 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C374 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C375 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C376 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C377 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C378 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C379 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C380 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C381 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C382 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C383 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C384 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C385 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C386 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.843945f
C387 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C388 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.49679f
C389 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C390 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C391 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C392 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C393 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C394 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C395 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C396 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C397 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.425359f
C398 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 34.661938f
C399 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C400 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C401 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C402 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C403 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C404 cp2_buffer_5stage_0/cp2_buffer1_1/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.270148f
C405 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C406 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.234749f
C407 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C408 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C409 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C410 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C411 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C412 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C413 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C414 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C415 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C416 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C417 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C418 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C419 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C420 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C421 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C422 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.064581f
C423 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C424 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.91548f
C425 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C426 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C427 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C428 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C429 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C430 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C431 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C432 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C433 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C434 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C435 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C436 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C437 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C438 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C439 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C440 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C441 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C442 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C443 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C444 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C445 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C446 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C447 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C448 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 49.246037f
C449 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.843945f
C450 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C451 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.49679f
C452 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C453 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C454 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C455 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C456 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C457 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C458 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C459 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C460 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.425359f
C461 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.292723f
C462 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C463 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C464 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C465 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C466 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C467 cp2_buffer_5stage_0/cp2_buffer1_2/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.081805f
C468 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C469 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C470 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C471 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C472 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C473 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C474 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C475 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C476 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C477 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C478 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C479 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C480 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C481 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C482 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C483 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C484 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C485 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.031953f
C486 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C487 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.29302f
C488 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C489 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C490 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C491 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C492 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C493 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C494 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C495 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C496 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C497 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C498 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C499 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C500 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C501 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C502 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C503 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C504 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C505 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C506 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C507 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C508 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C509 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C510 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C511 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C512 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C513 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.95876f
C514 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C515 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C516 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C517 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C518 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C519 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C520 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C521 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C522 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
C523 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 24.346807f
C524 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C525 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C526 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C527 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C528 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C529 cp2_buffer_5stage_0/cp2_buffer2_1/buffer_digital_2/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.84415f
C530 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C531 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C532 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C533 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C534 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C535 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C536 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C537 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C538 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C539 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C540 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C541 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C542 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C543 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C544 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in7 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 50.792114f
C545 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C546 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C547 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C548 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.031953f
C549 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C550 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.29452f
C551 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C552 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C553 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C554 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C555 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C556 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C557 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C558 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C559 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C560 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C561 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C562 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C563 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C564 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C565 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C566 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C567 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C568 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C569 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C570 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C571 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C572 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C573 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C574 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C575 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C576 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.97966f
C577 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C578 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C579 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C580 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C581 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C582 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C583 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C584 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C585 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
C586 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C587 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C588 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C589 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C590 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C591 cp2_buffer_5stage_0/cp2_buffer2_0/buffer_digital_2/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.985027f
C592 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C593 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43748f
C594 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C595 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C596 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C597 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C598 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C599 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C600 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/in5 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 36.018192f
C601 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C602 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C603 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C604 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C605 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C606 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C607 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C608 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C609 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C610 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.031953f
C611 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C612 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.29622f
C613 cp1_buffer_5stage_0/cp1_buffer1_2/vdd cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.81501p
C614 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C615 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C616 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C617 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C618 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C619 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C620 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C621 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C622 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C623 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C624 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C625 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C626 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C627 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C628 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C629 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C630 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C631 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C632 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C633 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C634 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C635 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C636 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C637 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.390842f
C638 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C639 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.97966f
C640 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C641 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C642 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C643 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C644 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C645 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C646 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C647 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.581652f
C648 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.634558f
C649 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.596436f
C650 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C651 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C652 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C653 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C654 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C655 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C656 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C657 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C658 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C659 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C660 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C661 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C662 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.33176f
C663 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.21436f
C664 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.683598f
C665 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C666 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C667 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C668 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C669 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C670 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C671 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C672 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C673 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C674 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C675 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C676 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C677 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C678 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C679 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C680 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C681 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C682 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C683 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C684 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C685 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C686 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C687 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C688 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C689 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C690 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C691 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C692 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C693 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C694 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C695 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C696 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 94.613235f
C697 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C698 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C699 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C700 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 0.10133p
C701 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C702 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C703 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C704 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C705 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C706 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C707 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C708 cp1_buffer_5stage_0/cp1_buffer1_2/clk_in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 5.346588f
C709 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C710 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.596436f
C711 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C712 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C713 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C714 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C715 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C716 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C717 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C718 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C719 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C720 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C721 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C722 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C723 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.33176f
C724 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.21436f
C725 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.683598f
C726 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C727 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C728 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C729 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C730 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C731 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C732 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C733 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C734 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C735 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C736 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C737 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C738 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C739 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C740 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C741 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C742 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C743 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C744 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C745 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C746 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C747 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C748 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C749 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C750 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C751 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C752 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C753 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C754 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C755 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C756 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C757 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 94.613235f
C758 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C759 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C760 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C761 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 0.10133p
C762 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C763 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C764 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C765 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C766 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C767 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C768 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C769 cp1_buffer_5stage_0/cp1_buffer1_1/clk_in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 4.427201f
C770 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C771 cp1_buffer_5stage_0/cp1_buffer1_2/clk_out cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.510713f
C772 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.463037f
C773 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.175129f
C774 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C775 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C776 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C777 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C778 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C779 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C780 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C781 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C782 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C783 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C784 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C785 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C786 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.771611f
C787 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.538747f
C788 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C789 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C790 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C791 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C792 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C793 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C794 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C795 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C796 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C797 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C798 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C799 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C800 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C801 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C802 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C803 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C804 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C805 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C806 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C807 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C808 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C809 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C810 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C811 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C812 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C813 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C814 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C815 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C816 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C817 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C818 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C819 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89.87499f
C820 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C821 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C822 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C823 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89.042244f
C824 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C825 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C826 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C827 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C828 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C829 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C830 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C831 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C832 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.344427f
C833 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 40.144115f
C834 cp1_buffer_5stage_0/cp1_buffer1_1/clk_out cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.469013f
C835 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.463037f
C836 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.175129f
C837 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C838 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C839 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C840 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C841 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C842 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C843 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C844 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C845 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C846 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C847 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C848 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C849 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.771611f
C850 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.538747f
C851 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.476783f
C852 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C853 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C854 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C855 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C856 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C857 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C858 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C859 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C860 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C861 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C862 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C863 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C864 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C865 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C866 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C867 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C868 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C869 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C870 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C871 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C872 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C873 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C874 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C875 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C876 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C877 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C878 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C879 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C880 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C881 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C882 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C883 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89.87499f
C884 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C885 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C886 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C887 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89.042244f
C888 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C889 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C890 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C891 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C892 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C893 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C894 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C895 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C896 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.344427f
C897 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 13.208359f
C898 cp1_buffer_5stage_0/cp1_buffer1_0/clk_in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 66.95308f
C899 cp1_buffer_5stage_0/cp1_buffer1_0/clk_out cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.485913f
C900 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.463037f
C901 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.175129f
C902 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C903 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C904 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C905 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C906 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C907 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C908 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C909 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C910 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C911 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C912 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C913 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C914 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.771611f
C915 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.538747f
C916 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.603806f
C917 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C918 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C919 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C920 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C921 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C922 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C923 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C924 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C925 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C926 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C927 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C928 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C929 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C930 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C931 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C932 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C933 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C934 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C935 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C936 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C937 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C938 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C939 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C940 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C941 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C942 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C943 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C944 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C945 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C946 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C947 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C948 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89.87499f
C949 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C950 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C951 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.337696f
C952 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89.01839f
C953 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.978376f
C954 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.608221f
C955 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C956 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C957 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.809951f
C958 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.172722f
C959 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.381627f
C960 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.834443f
C961 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.344427f
C962 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 10.368401f
.ends

