magic
tech sky130A
magscale 1 2
timestamp 1699130246
<< nwell >>
rect -1458 1760 -874 2212
rect 1358 2174 4094 2212
rect 1358 2156 4190 2174
rect 1426 2152 4190 2156
rect 1468 1760 4190 2152
<< nmos >>
rect 1566 1398 1596 1482
rect 1662 1398 1692 1482
rect 1758 1398 1788 1482
rect 1854 1398 1884 1482
rect 1950 1398 1980 1482
rect 2046 1398 2076 1482
rect 2142 1398 2172 1482
rect 2238 1398 2268 1482
rect 2334 1398 2364 1482
rect 2430 1398 2460 1482
rect 2526 1398 2556 1482
rect 2622 1398 2652 1482
rect 2718 1398 2748 1482
rect 2814 1398 2844 1482
rect 2910 1398 2940 1482
rect 3006 1398 3036 1482
rect 3102 1398 3132 1482
rect 3198 1398 3228 1482
rect 3294 1398 3324 1482
rect 3390 1398 3420 1482
rect 3486 1398 3516 1482
rect 3582 1398 3612 1482
rect 3678 1398 3708 1482
rect 3774 1398 3804 1482
rect 3870 1398 3900 1482
rect 3966 1398 3996 1482
rect 4062 1398 4092 1482
<< pmos >>
rect 1566 1860 1596 2112
rect 1662 1860 1692 2112
rect 1758 1860 1788 2112
rect 1854 1860 1884 2112
rect 1950 1860 1980 2112
rect 2046 1860 2076 2112
rect 2142 1860 2172 2112
rect 2238 1860 2268 2112
rect 2334 1860 2364 2112
rect 2430 1860 2460 2112
rect 2526 1860 2556 2112
rect 2622 1860 2652 2112
rect 2718 1860 2748 2112
rect 2814 1860 2844 2112
rect 2910 1860 2940 2112
rect 3006 1860 3036 2112
rect 3102 1860 3132 2112
rect 3198 1860 3228 2112
rect 3294 1860 3324 2112
rect 3390 1860 3420 2112
rect 3486 1860 3516 2112
rect 3582 1860 3612 2112
rect 3678 1860 3708 2112
rect 3774 1860 3804 2112
rect 3870 1860 3900 2112
rect 3966 1860 3996 2112
rect 4062 1860 4092 2112
<< ndiff >>
rect 1504 1470 1566 1482
rect 1504 1410 1516 1470
rect 1550 1410 1566 1470
rect 1504 1398 1566 1410
rect 1596 1470 1662 1482
rect 1596 1410 1612 1470
rect 1646 1410 1662 1470
rect 1596 1398 1662 1410
rect 1692 1470 1758 1482
rect 1692 1410 1708 1470
rect 1742 1410 1758 1470
rect 1692 1398 1758 1410
rect 1788 1470 1854 1482
rect 1788 1410 1804 1470
rect 1838 1410 1854 1470
rect 1788 1398 1854 1410
rect 1884 1470 1950 1482
rect 1884 1410 1900 1470
rect 1934 1410 1950 1470
rect 1884 1398 1950 1410
rect 1980 1470 2046 1482
rect 1980 1410 1996 1470
rect 2030 1410 2046 1470
rect 1980 1398 2046 1410
rect 2076 1470 2142 1482
rect 2076 1410 2092 1470
rect 2126 1410 2142 1470
rect 2076 1398 2142 1410
rect 2172 1470 2238 1482
rect 2172 1410 2188 1470
rect 2222 1410 2238 1470
rect 2172 1398 2238 1410
rect 2268 1470 2334 1482
rect 2268 1410 2284 1470
rect 2318 1410 2334 1470
rect 2268 1398 2334 1410
rect 2364 1470 2430 1482
rect 2364 1410 2380 1470
rect 2414 1410 2430 1470
rect 2364 1398 2430 1410
rect 2460 1470 2526 1482
rect 2460 1410 2476 1470
rect 2510 1410 2526 1470
rect 2460 1398 2526 1410
rect 2556 1470 2622 1482
rect 2556 1410 2572 1470
rect 2606 1410 2622 1470
rect 2556 1398 2622 1410
rect 2652 1470 2718 1482
rect 2652 1410 2668 1470
rect 2702 1410 2718 1470
rect 2652 1398 2718 1410
rect 2748 1470 2814 1482
rect 2748 1410 2764 1470
rect 2798 1410 2814 1470
rect 2748 1398 2814 1410
rect 2844 1470 2910 1482
rect 2844 1410 2860 1470
rect 2894 1410 2910 1470
rect 2844 1398 2910 1410
rect 2940 1470 3006 1482
rect 2940 1410 2956 1470
rect 2990 1410 3006 1470
rect 2940 1398 3006 1410
rect 3036 1470 3102 1482
rect 3036 1410 3052 1470
rect 3086 1410 3102 1470
rect 3036 1398 3102 1410
rect 3132 1470 3198 1482
rect 3132 1410 3148 1470
rect 3182 1410 3198 1470
rect 3132 1398 3198 1410
rect 3228 1470 3294 1482
rect 3228 1410 3244 1470
rect 3278 1410 3294 1470
rect 3228 1398 3294 1410
rect 3324 1470 3390 1482
rect 3324 1410 3340 1470
rect 3374 1410 3390 1470
rect 3324 1398 3390 1410
rect 3420 1470 3486 1482
rect 3420 1410 3436 1470
rect 3470 1410 3486 1470
rect 3420 1398 3486 1410
rect 3516 1470 3582 1482
rect 3516 1410 3532 1470
rect 3566 1410 3582 1470
rect 3516 1398 3582 1410
rect 3612 1470 3678 1482
rect 3612 1410 3628 1470
rect 3662 1410 3678 1470
rect 3612 1398 3678 1410
rect 3708 1470 3774 1482
rect 3708 1410 3724 1470
rect 3758 1410 3774 1470
rect 3708 1398 3774 1410
rect 3804 1470 3870 1482
rect 3804 1410 3820 1470
rect 3854 1410 3870 1470
rect 3804 1398 3870 1410
rect 3900 1470 3966 1482
rect 3900 1410 3916 1470
rect 3950 1410 3966 1470
rect 3900 1398 3966 1410
rect 3996 1470 4062 1482
rect 3996 1410 4012 1470
rect 4046 1410 4062 1470
rect 3996 1398 4062 1410
rect 4092 1470 4154 1482
rect 4092 1410 4108 1470
rect 4142 1410 4154 1470
rect 4092 1398 4154 1410
<< pdiff >>
rect 1504 2100 1566 2112
rect 1504 1872 1516 2100
rect 1550 1872 1566 2100
rect 1504 1860 1566 1872
rect 1596 2100 1662 2112
rect 1596 1872 1612 2100
rect 1646 1872 1662 2100
rect 1596 1860 1662 1872
rect 1692 2100 1758 2112
rect 1692 1872 1708 2100
rect 1742 1872 1758 2100
rect 1692 1860 1758 1872
rect 1788 2100 1854 2112
rect 1788 1872 1804 2100
rect 1838 1872 1854 2100
rect 1788 1860 1854 1872
rect 1884 2100 1950 2112
rect 1884 1872 1900 2100
rect 1934 1872 1950 2100
rect 1884 1860 1950 1872
rect 1980 2100 2046 2112
rect 1980 1872 1996 2100
rect 2030 1872 2046 2100
rect 1980 1860 2046 1872
rect 2076 2100 2142 2112
rect 2076 1872 2092 2100
rect 2126 1872 2142 2100
rect 2076 1860 2142 1872
rect 2172 2100 2238 2112
rect 2172 1872 2188 2100
rect 2222 1872 2238 2100
rect 2172 1860 2238 1872
rect 2268 2100 2334 2112
rect 2268 1872 2284 2100
rect 2318 1872 2334 2100
rect 2268 1860 2334 1872
rect 2364 2100 2430 2112
rect 2364 1872 2380 2100
rect 2414 1872 2430 2100
rect 2364 1860 2430 1872
rect 2460 2100 2526 2112
rect 2460 1872 2476 2100
rect 2510 1872 2526 2100
rect 2460 1860 2526 1872
rect 2556 2100 2622 2112
rect 2556 1872 2572 2100
rect 2606 1872 2622 2100
rect 2556 1860 2622 1872
rect 2652 2100 2718 2112
rect 2652 1872 2668 2100
rect 2702 1872 2718 2100
rect 2652 1860 2718 1872
rect 2748 2100 2814 2112
rect 2748 1872 2764 2100
rect 2798 1872 2814 2100
rect 2748 1860 2814 1872
rect 2844 2100 2910 2112
rect 2844 1872 2860 2100
rect 2894 1872 2910 2100
rect 2844 1860 2910 1872
rect 2940 2100 3006 2112
rect 2940 1872 2956 2100
rect 2990 1872 3006 2100
rect 2940 1860 3006 1872
rect 3036 2100 3102 2112
rect 3036 1872 3052 2100
rect 3086 1872 3102 2100
rect 3036 1860 3102 1872
rect 3132 2100 3198 2112
rect 3132 1872 3148 2100
rect 3182 1872 3198 2100
rect 3132 1860 3198 1872
rect 3228 2100 3294 2112
rect 3228 1872 3244 2100
rect 3278 1872 3294 2100
rect 3228 1860 3294 1872
rect 3324 2100 3390 2112
rect 3324 1872 3340 2100
rect 3374 1872 3390 2100
rect 3324 1860 3390 1872
rect 3420 2100 3486 2112
rect 3420 1872 3436 2100
rect 3470 1872 3486 2100
rect 3420 1860 3486 1872
rect 3516 2100 3582 2112
rect 3516 1872 3532 2100
rect 3566 1872 3582 2100
rect 3516 1860 3582 1872
rect 3612 2100 3678 2112
rect 3612 1872 3628 2100
rect 3662 1872 3678 2100
rect 3612 1860 3678 1872
rect 3708 2100 3774 2112
rect 3708 1872 3724 2100
rect 3758 1872 3774 2100
rect 3708 1860 3774 1872
rect 3804 2100 3870 2112
rect 3804 1872 3820 2100
rect 3854 1872 3870 2100
rect 3804 1860 3870 1872
rect 3900 2100 3966 2112
rect 3900 1872 3916 2100
rect 3950 1872 3966 2100
rect 3900 1860 3966 1872
rect 3996 2100 4062 2112
rect 3996 1872 4012 2100
rect 4046 1872 4062 2100
rect 3996 1860 4062 1872
rect 4092 2100 4154 2112
rect 4092 1872 4108 2100
rect 4142 1872 4154 2100
rect 4092 1860 4154 1872
<< ndiffc >>
rect 1516 1410 1550 1470
rect 1612 1410 1646 1470
rect 1708 1410 1742 1470
rect 1804 1410 1838 1470
rect 1900 1410 1934 1470
rect 1996 1410 2030 1470
rect 2092 1410 2126 1470
rect 2188 1410 2222 1470
rect 2284 1410 2318 1470
rect 2380 1410 2414 1470
rect 2476 1410 2510 1470
rect 2572 1410 2606 1470
rect 2668 1410 2702 1470
rect 2764 1410 2798 1470
rect 2860 1410 2894 1470
rect 2956 1410 2990 1470
rect 3052 1410 3086 1470
rect 3148 1410 3182 1470
rect 3244 1410 3278 1470
rect 3340 1410 3374 1470
rect 3436 1410 3470 1470
rect 3532 1410 3566 1470
rect 3628 1410 3662 1470
rect 3724 1410 3758 1470
rect 3820 1410 3854 1470
rect 3916 1410 3950 1470
rect 4012 1410 4046 1470
rect 4108 1410 4142 1470
<< pdiffc >>
rect 1516 1872 1550 2100
rect 1612 1872 1646 2100
rect 1708 1872 1742 2100
rect 1804 1872 1838 2100
rect 1900 1872 1934 2100
rect 1996 1872 2030 2100
rect 2092 1872 2126 2100
rect 2188 1872 2222 2100
rect 2284 1872 2318 2100
rect 2380 1872 2414 2100
rect 2476 1872 2510 2100
rect 2572 1872 2606 2100
rect 2668 1872 2702 2100
rect 2764 1872 2798 2100
rect 2860 1872 2894 2100
rect 2956 1872 2990 2100
rect 3052 1872 3086 2100
rect 3148 1872 3182 2100
rect 3244 1872 3278 2100
rect 3340 1872 3374 2100
rect 3436 1872 3470 2100
rect 3532 1872 3566 2100
rect 3628 1872 3662 2100
rect 3724 1872 3758 2100
rect 3820 1872 3854 2100
rect 3916 1872 3950 2100
rect 4012 1872 4046 2100
rect 4108 1872 4142 2100
<< psubdiff >>
rect -1354 1456 -1262 1482
rect -1354 1392 -1336 1456
rect -1280 1392 -1262 1456
rect -1354 1366 -1262 1392
<< nsubdiff >>
rect -1378 2124 -1292 2166
rect -1378 1978 -1356 2124
rect -1312 1978 -1292 2124
rect -1378 1938 -1292 1978
<< psubdiffcont >>
rect -1336 1392 -1280 1456
<< nsubdiffcont >>
rect -1356 1978 -1312 2124
<< poly >>
rect 206 2194 236 2198
rect 1644 2194 1710 2209
rect 1836 2194 1902 2209
rect 2028 2194 2094 2209
rect 2220 2194 2286 2209
rect 2412 2194 2478 2209
rect 2604 2194 2670 2209
rect 2796 2194 2862 2209
rect 2910 2194 2940 2198
rect 2988 2194 3054 2209
rect 3180 2194 3246 2209
rect 3372 2194 3438 2209
rect 3564 2194 3630 2209
rect 3756 2194 3822 2209
rect 3948 2194 4014 2209
rect -1140 2162 1390 2194
rect 1564 2193 4094 2194
rect 1564 2162 1660 2193
rect -1138 2114 -1108 2162
rect -946 2114 -916 2162
rect -754 2114 -724 2162
rect -562 2116 -532 2162
rect -370 2114 -340 2162
rect -178 2118 -148 2162
rect 14 2116 44 2162
rect 206 2122 236 2162
rect 398 2114 428 2162
rect 590 2118 620 2162
rect 782 2118 812 2162
rect 974 2118 1004 2162
rect 1166 2118 1196 2162
rect 1358 2116 1388 2162
rect 1566 2112 1596 2162
rect 1644 2159 1660 2162
rect 1694 2162 1852 2193
rect 1694 2159 1710 2162
rect 1644 2143 1710 2159
rect 1662 2112 1692 2143
rect 1758 2112 1788 2162
rect 1836 2159 1852 2162
rect 1886 2162 2044 2193
rect 1886 2159 1902 2162
rect 1836 2143 1902 2159
rect 1854 2112 1884 2143
rect 1950 2112 1980 2162
rect 2028 2159 2044 2162
rect 2078 2162 2236 2193
rect 2078 2159 2094 2162
rect 2028 2143 2094 2159
rect 2046 2112 2076 2143
rect 2142 2112 2172 2162
rect 2220 2159 2236 2162
rect 2270 2162 2428 2193
rect 2270 2159 2286 2162
rect 2220 2143 2286 2159
rect 2238 2112 2268 2143
rect 2334 2112 2364 2162
rect 2412 2159 2428 2162
rect 2462 2162 2620 2193
rect 2462 2159 2478 2162
rect 2412 2143 2478 2159
rect 2430 2112 2460 2143
rect 2526 2112 2556 2162
rect 2604 2159 2620 2162
rect 2654 2162 2812 2193
rect 2654 2159 2670 2162
rect 2604 2143 2670 2159
rect 2622 2112 2652 2143
rect 2718 2112 2748 2162
rect 2796 2159 2812 2162
rect 2846 2162 3004 2193
rect 2846 2159 2862 2162
rect 2796 2143 2862 2159
rect 2814 2112 2844 2143
rect 2910 2112 2940 2162
rect 2988 2159 3004 2162
rect 3038 2162 3196 2193
rect 3038 2159 3054 2162
rect 2988 2143 3054 2159
rect 3006 2112 3036 2143
rect 3102 2112 3132 2162
rect 3180 2159 3196 2162
rect 3230 2162 3388 2193
rect 3230 2159 3246 2162
rect 3180 2143 3246 2159
rect 3198 2112 3228 2143
rect 3294 2112 3324 2162
rect 3372 2159 3388 2162
rect 3422 2162 3580 2193
rect 3422 2159 3438 2162
rect 3372 2143 3438 2159
rect 3390 2112 3420 2143
rect 3486 2112 3516 2162
rect 3564 2159 3580 2162
rect 3614 2162 3772 2193
rect 3614 2159 3630 2162
rect 3564 2143 3630 2159
rect 3582 2112 3612 2143
rect 3678 2112 3708 2162
rect 3756 2159 3772 2162
rect 3806 2162 3964 2193
rect 3806 2159 3822 2162
rect 3756 2143 3822 2159
rect 3774 2112 3804 2143
rect 3870 2112 3900 2162
rect 3948 2159 3964 2162
rect 3998 2162 4094 2193
rect 3998 2159 4014 2162
rect 3948 2143 4014 2159
rect 3966 2112 3996 2143
rect 4062 2112 4092 2162
rect -1138 1812 -1108 1845
rect -1042 1812 -1012 1856
rect -850 1812 -820 1856
rect -658 1812 -628 1856
rect -466 1812 -436 1856
rect -274 1812 -244 1858
rect -82 1812 -52 1856
rect 110 1812 140 1856
rect 302 1812 332 1858
rect 494 1812 524 1856
rect 686 1812 716 1858
rect 878 1812 908 1856
rect 1070 1812 1100 1856
rect 1262 1812 1292 1856
rect 1566 1829 1596 1860
rect 1548 1813 1614 1829
rect 1548 1812 1564 1813
rect -1158 1778 1391 1812
rect 1546 1779 1564 1812
rect 1598 1812 1614 1813
rect 1662 1812 1692 1860
rect 1758 1829 1788 1860
rect 1740 1813 1806 1829
rect 1740 1812 1756 1813
rect 1598 1779 1756 1812
rect 1790 1812 1806 1813
rect 1854 1812 1884 1860
rect 1950 1829 1980 1860
rect 1932 1813 1998 1829
rect 1932 1812 1948 1813
rect 1790 1779 1948 1812
rect 1982 1812 1998 1813
rect 2046 1812 2076 1860
rect 2142 1829 2172 1860
rect 2124 1813 2190 1829
rect 2124 1812 2140 1813
rect 1982 1779 2140 1812
rect 2174 1812 2190 1813
rect 2238 1812 2268 1860
rect 2334 1829 2364 1860
rect 2316 1813 2382 1829
rect 2316 1812 2332 1813
rect 2174 1779 2332 1812
rect 2366 1812 2382 1813
rect 2430 1812 2460 1860
rect 2526 1829 2556 1860
rect 2508 1813 2574 1829
rect 2508 1812 2524 1813
rect 2366 1779 2524 1812
rect 2558 1812 2574 1813
rect 2622 1812 2652 1860
rect 2718 1829 2748 1860
rect 2700 1813 2766 1829
rect 2700 1812 2716 1813
rect 2558 1779 2716 1812
rect 2750 1812 2766 1813
rect 2814 1812 2844 1860
rect 2910 1829 2940 1860
rect 2892 1813 2958 1829
rect 2892 1812 2908 1813
rect 2750 1779 2908 1812
rect 2942 1812 2958 1813
rect 3006 1812 3036 1860
rect 3102 1829 3132 1860
rect 3084 1813 3150 1829
rect 3084 1812 3100 1813
rect 2942 1779 3100 1812
rect 3134 1812 3150 1813
rect 3198 1812 3228 1860
rect 3294 1829 3324 1860
rect 3276 1813 3342 1829
rect 3276 1812 3292 1813
rect 3134 1779 3292 1812
rect 3326 1812 3342 1813
rect 3390 1812 3420 1860
rect 3486 1829 3516 1860
rect 3468 1813 3534 1829
rect 3468 1812 3484 1813
rect 3326 1779 3484 1812
rect 3518 1812 3534 1813
rect 3582 1812 3612 1860
rect 3678 1829 3708 1860
rect 3660 1813 3726 1829
rect 3660 1812 3676 1813
rect 3518 1779 3676 1812
rect 3710 1812 3726 1813
rect 3774 1812 3804 1860
rect 3870 1829 3900 1860
rect 3852 1813 3918 1829
rect 3852 1812 3868 1813
rect 3710 1779 3868 1812
rect 3902 1812 3918 1813
rect 3966 1812 3996 1860
rect 4062 1829 4092 1860
rect 4044 1813 4110 1829
rect 4044 1812 4060 1813
rect 3902 1779 4060 1812
rect 4094 1779 4110 1813
rect 1546 1778 4110 1779
rect -1138 1555 -1108 1778
rect -562 1555 -532 1556
rect 974 1555 1004 1556
rect 1166 1555 1196 1556
rect 1357 1555 1391 1778
rect 1548 1763 1614 1778
rect 1740 1763 1806 1778
rect 1932 1763 1998 1778
rect 2124 1763 2190 1778
rect 2316 1763 2382 1778
rect 2508 1763 2574 1778
rect 2700 1763 2766 1778
rect 2892 1763 2958 1778
rect 3084 1763 3150 1778
rect 3276 1763 3342 1778
rect 3468 1763 3534 1778
rect 3660 1763 3726 1778
rect 3852 1763 3918 1778
rect 4044 1763 4110 1778
rect 1566 1680 1596 1763
rect -1139 1521 1391 1555
rect 1436 1666 1598 1680
rect 1436 1564 1454 1666
rect 1582 1564 1598 1666
rect 1436 1556 1598 1564
rect 1644 1556 1710 1570
rect 1436 1555 1710 1556
rect 1836 1555 1902 1570
rect 2028 1555 2094 1570
rect 2142 1555 2172 1556
rect 2220 1555 2286 1570
rect 2412 1555 2478 1570
rect 2604 1555 2670 1570
rect 2796 1555 2862 1570
rect 2988 1555 3054 1570
rect 3180 1555 3246 1570
rect 3372 1555 3438 1570
rect 3564 1555 3630 1570
rect 3678 1555 3708 1556
rect 3756 1555 3822 1570
rect 3870 1555 3900 1556
rect 3948 1555 4014 1570
rect 4061 1555 4095 1763
rect 1436 1554 4095 1555
rect 1436 1552 1660 1554
rect 1565 1521 1660 1552
rect -1138 1482 -1108 1521
rect -946 1484 -916 1521
rect -754 1486 -724 1521
rect -562 1488 -532 1521
rect -370 1486 -340 1521
rect -178 1486 -148 1521
rect 14 1486 44 1521
rect 206 1486 236 1521
rect 398 1486 428 1521
rect 590 1486 620 1521
rect 782 1484 812 1521
rect 974 1488 1004 1521
rect 1166 1488 1196 1521
rect 1358 1488 1388 1521
rect 1566 1520 1660 1521
rect 1694 1521 1852 1554
rect 1694 1520 1710 1521
rect 1566 1482 1596 1520
rect 1644 1504 1710 1520
rect 1662 1482 1692 1504
rect 1758 1482 1788 1521
rect 1836 1520 1852 1521
rect 1886 1521 2044 1554
rect 1886 1520 1902 1521
rect 1836 1504 1902 1520
rect 1854 1482 1884 1504
rect 1950 1482 1980 1521
rect 2028 1520 2044 1521
rect 2078 1521 2236 1554
rect 2078 1520 2094 1521
rect 2028 1504 2094 1520
rect 2046 1482 2076 1504
rect 2142 1482 2172 1521
rect 2220 1520 2236 1521
rect 2270 1521 2428 1554
rect 2270 1520 2286 1521
rect 2220 1504 2286 1520
rect 2238 1482 2268 1504
rect 2334 1482 2364 1521
rect 2412 1520 2428 1521
rect 2462 1521 2620 1554
rect 2462 1520 2478 1521
rect 2412 1504 2478 1520
rect 2430 1482 2460 1504
rect 2526 1482 2556 1521
rect 2604 1520 2620 1521
rect 2654 1521 2812 1554
rect 2654 1520 2670 1521
rect 2604 1504 2670 1520
rect 2622 1482 2652 1504
rect 2718 1482 2748 1521
rect 2796 1520 2812 1521
rect 2846 1521 3004 1554
rect 2846 1520 2862 1521
rect 2796 1504 2862 1520
rect 2814 1482 2844 1504
rect 2910 1482 2940 1521
rect 2988 1520 3004 1521
rect 3038 1521 3196 1554
rect 3038 1520 3054 1521
rect 2988 1504 3054 1520
rect 3006 1482 3036 1504
rect 3102 1482 3132 1521
rect 3180 1520 3196 1521
rect 3230 1521 3388 1554
rect 3230 1520 3246 1521
rect 3180 1504 3246 1520
rect 3198 1482 3228 1504
rect 3294 1482 3324 1521
rect 3372 1520 3388 1521
rect 3422 1521 3580 1554
rect 3422 1520 3438 1521
rect 3372 1504 3438 1520
rect 3390 1482 3420 1504
rect 3486 1482 3516 1521
rect 3564 1520 3580 1521
rect 3614 1521 3772 1554
rect 3614 1520 3630 1521
rect 3564 1504 3630 1520
rect 3582 1482 3612 1504
rect 3678 1482 3708 1521
rect 3756 1520 3772 1521
rect 3806 1521 3964 1554
rect 3806 1520 3822 1521
rect 3756 1504 3822 1520
rect 3774 1482 3804 1504
rect 3870 1482 3900 1521
rect 3948 1520 3964 1521
rect 3998 1521 4095 1554
rect 3998 1520 4014 1521
rect 3948 1504 4014 1520
rect 3966 1482 3996 1504
rect 4062 1482 4092 1521
rect -1042 1360 -1012 1398
rect -850 1360 -820 1398
rect -658 1360 -628 1398
rect -466 1360 -436 1408
rect -274 1360 -244 1398
rect -82 1360 -52 1396
rect 110 1360 140 1394
rect 302 1360 332 1394
rect 494 1360 524 1394
rect 686 1360 716 1394
rect 878 1360 908 1398
rect 1070 1360 1100 1394
rect 1262 1360 1292 1396
rect 1566 1376 1596 1398
rect 1548 1360 1614 1376
rect 1662 1360 1692 1398
rect 1758 1376 1788 1398
rect 1740 1360 1806 1376
rect 1854 1360 1884 1398
rect 1950 1376 1980 1398
rect 1932 1360 1998 1376
rect 2046 1360 2076 1398
rect 2142 1376 2172 1398
rect 2124 1360 2190 1376
rect 2238 1360 2268 1398
rect 2334 1376 2364 1398
rect 2316 1360 2382 1376
rect 2430 1360 2460 1398
rect 2526 1376 2556 1398
rect 2508 1360 2574 1376
rect 2622 1360 2652 1398
rect 2718 1376 2748 1398
rect 2700 1360 2766 1376
rect 2814 1360 2844 1398
rect 2910 1376 2940 1398
rect 2892 1360 2958 1376
rect 3006 1360 3036 1398
rect 3102 1376 3132 1398
rect 3084 1360 3150 1376
rect 3198 1360 3228 1398
rect 3294 1376 3324 1398
rect 3276 1360 3342 1376
rect 3390 1360 3420 1398
rect 3486 1376 3516 1398
rect 3468 1360 3534 1376
rect 3582 1360 3612 1398
rect 3678 1376 3708 1398
rect 3660 1360 3726 1376
rect 3774 1360 3804 1398
rect 3870 1376 3900 1398
rect 3852 1360 3918 1376
rect 3966 1360 3996 1398
rect 4062 1376 4092 1398
rect 4044 1360 4110 1376
rect -1157 1326 1406 1360
rect 1547 1326 1564 1360
rect 1598 1326 1756 1360
rect 1790 1326 1948 1360
rect 1982 1326 2140 1360
rect 2174 1326 2332 1360
rect 2366 1326 2524 1360
rect 2558 1326 2716 1360
rect 2750 1326 2908 1360
rect 2942 1326 3100 1360
rect 3134 1326 3292 1360
rect 3326 1326 3484 1360
rect 3518 1326 3676 1360
rect 3710 1326 3868 1360
rect 3902 1326 4060 1360
rect 4094 1326 4110 1360
rect 1548 1310 1614 1326
rect 1740 1310 1806 1326
rect 1932 1310 1998 1326
rect 2124 1310 2190 1326
rect 2316 1310 2382 1326
rect 2508 1310 2574 1326
rect 2700 1310 2766 1326
rect 2892 1310 2958 1326
rect 3084 1310 3150 1326
rect 3276 1310 3342 1326
rect 3468 1310 3534 1326
rect 3660 1310 3726 1326
rect 3852 1310 3918 1326
rect 4044 1310 4110 1326
<< polycont >>
rect 1660 2159 1694 2193
rect 1852 2159 1886 2193
rect 2044 2159 2078 2193
rect 2236 2159 2270 2193
rect 2428 2159 2462 2193
rect 2620 2159 2654 2193
rect 2812 2159 2846 2193
rect 3004 2159 3038 2193
rect 3196 2159 3230 2193
rect 3388 2159 3422 2193
rect 3580 2159 3614 2193
rect 3772 2159 3806 2193
rect 3964 2159 3998 2193
rect 1564 1779 1598 1813
rect 1756 1779 1790 1813
rect 1948 1779 1982 1813
rect 2140 1779 2174 1813
rect 2332 1779 2366 1813
rect 2524 1779 2558 1813
rect 2716 1779 2750 1813
rect 2908 1779 2942 1813
rect 3100 1779 3134 1813
rect 3292 1779 3326 1813
rect 3484 1779 3518 1813
rect 3676 1779 3710 1813
rect 3868 1779 3902 1813
rect 4060 1779 4094 1813
rect 1454 1564 1582 1666
rect 1660 1520 1694 1554
rect 1852 1520 1886 1554
rect 2044 1520 2078 1554
rect 2236 1520 2270 1554
rect 2428 1520 2462 1554
rect 2620 1520 2654 1554
rect 2812 1520 2846 1554
rect 3004 1520 3038 1554
rect 3196 1520 3230 1554
rect 3388 1520 3422 1554
rect 3580 1520 3614 1554
rect 3772 1520 3806 1554
rect 3964 1520 3998 1554
rect 1564 1326 1598 1360
rect 1756 1326 1790 1360
rect 1948 1326 1982 1360
rect 2140 1326 2174 1360
rect 2332 1326 2366 1360
rect 2524 1326 2558 1360
rect 2716 1326 2750 1360
rect 2908 1326 2942 1360
rect 3100 1326 3134 1360
rect 3292 1326 3326 1360
rect 3484 1326 3518 1360
rect 3676 1326 3710 1360
rect 3868 1326 3902 1360
rect 4060 1326 4094 1360
<< locali >>
rect -1061 2192 1390 2194
rect 1643 2193 4094 2194
rect 1643 2192 1660 2193
rect -1378 2124 -1292 2166
rect -1140 2160 1390 2192
rect -1140 2158 -1044 2160
rect 1228 2158 1310 2160
rect 1564 2158 1660 2192
rect 1694 2160 1852 2193
rect 1694 2159 1710 2160
rect 1836 2159 1852 2160
rect 1886 2160 2044 2193
rect 1886 2159 1902 2160
rect 2028 2159 2044 2160
rect 2078 2160 2236 2193
rect 2078 2159 2094 2160
rect 2220 2159 2236 2160
rect 2270 2160 2428 2193
rect 2270 2159 2286 2160
rect 2412 2159 2428 2160
rect 2462 2160 2620 2193
rect 2462 2159 2478 2160
rect 2604 2159 2620 2160
rect 2654 2160 2812 2193
rect 2654 2159 2670 2160
rect 2796 2159 2812 2160
rect 2846 2160 3004 2193
rect 2846 2159 2862 2160
rect 2988 2159 3004 2160
rect 3038 2160 3196 2193
rect 3038 2159 3054 2160
rect 3180 2159 3196 2160
rect 3230 2160 3388 2193
rect 3230 2159 3246 2160
rect 3372 2159 3388 2160
rect 3422 2160 3580 2193
rect 3422 2159 3438 2160
rect 3564 2159 3580 2160
rect 3614 2160 3772 2193
rect 3614 2159 3630 2160
rect 3756 2159 3772 2160
rect 3806 2160 3964 2193
rect 3806 2159 3822 2160
rect 3932 2159 3964 2160
rect 3998 2160 4094 2193
rect 3998 2159 4014 2160
rect 3932 2158 4014 2159
rect -1378 1978 -1356 2124
rect -1312 1978 -1292 2124
rect -1378 1938 -1292 1978
rect 1516 2100 1550 2116
rect 1516 1856 1550 1872
rect 1612 2100 1646 2116
rect 1612 1856 1646 1872
rect 1708 2100 1742 2116
rect 1708 1856 1742 1872
rect 1804 2100 1838 2116
rect 1804 1856 1838 1872
rect 1900 2100 1934 2116
rect 1900 1856 1934 1872
rect 1996 2100 2030 2116
rect 1996 1856 2030 1872
rect 2092 2100 2126 2116
rect 2092 1856 2126 1872
rect 2188 2100 2222 2116
rect 2188 1856 2222 1872
rect 2284 2100 2318 2116
rect 2284 1856 2318 1872
rect 2380 2100 2414 2116
rect 2380 1856 2414 1872
rect 2476 2100 2510 2116
rect 2476 1856 2510 1872
rect 2572 2100 2606 2116
rect 2572 1856 2606 1872
rect 2668 2100 2702 2116
rect 2668 1856 2702 1872
rect 2764 2100 2798 2116
rect 2764 1856 2798 1872
rect 2860 2100 2894 2116
rect 2860 1856 2894 1872
rect 2956 2100 2990 2116
rect 2956 1856 2990 1872
rect 3052 2100 3086 2116
rect 3052 1856 3086 1872
rect 3148 2100 3182 2116
rect 3148 1856 3182 1872
rect 3244 2100 3278 2116
rect 3244 1856 3278 1872
rect 3340 2100 3374 2116
rect 3340 1856 3374 1872
rect 3436 2100 3470 2116
rect 3436 1856 3470 1872
rect 3532 2100 3566 2116
rect 3532 1856 3566 1872
rect 3628 2100 3662 2116
rect 3628 1856 3662 1872
rect 3724 2100 3758 2116
rect 3724 1856 3758 1872
rect 3820 2100 3854 2116
rect 3820 1856 3854 1872
rect 3916 2100 3950 2116
rect 3916 1856 3950 1872
rect 4012 2100 4046 2116
rect 4012 1856 4046 1872
rect 4108 2100 4142 2116
rect 4108 1856 4142 1872
rect -1156 1778 1390 1814
rect 1548 1813 4094 1814
rect 1548 1779 1564 1813
rect 1598 1779 1756 1813
rect 1790 1779 1948 1813
rect 1982 1779 2140 1813
rect 2174 1779 2332 1813
rect 2366 1779 2524 1813
rect 2558 1779 2716 1813
rect 2750 1779 2908 1813
rect 2942 1779 3100 1813
rect 3134 1779 3292 1813
rect 3326 1779 3484 1813
rect 3518 1779 3676 1813
rect 3710 1779 3868 1813
rect 3902 1779 4060 1813
rect 4094 1779 4110 1813
rect 1548 1778 4094 1779
rect 1354 1556 1390 1778
rect -1138 1520 1390 1556
rect 1430 1666 1604 1680
rect 1430 1564 1454 1666
rect 1582 1564 1604 1666
rect 1430 1556 1604 1564
rect 4058 1556 4094 1778
rect 1430 1554 4094 1556
rect 1430 1552 1660 1554
rect 1566 1520 1660 1552
rect 1694 1520 1852 1554
rect 1886 1520 2044 1554
rect 2078 1520 2236 1554
rect 2270 1520 2428 1554
rect 2462 1520 2620 1554
rect 2654 1520 2812 1554
rect 2846 1520 3004 1554
rect 3038 1520 3196 1554
rect 3230 1520 3388 1554
rect 3422 1520 3580 1554
rect 3614 1520 3772 1554
rect 3806 1520 3964 1554
rect 3998 1520 4094 1554
rect -1354 1456 -1262 1482
rect -1354 1392 -1336 1456
rect -1280 1392 -1262 1456
rect 1516 1470 1550 1486
rect 1516 1394 1550 1410
rect 1612 1470 1646 1486
rect 1612 1394 1646 1410
rect 1708 1470 1742 1486
rect 1708 1394 1742 1410
rect 1804 1470 1838 1486
rect 1804 1394 1838 1410
rect 1900 1470 1934 1486
rect 1900 1394 1934 1410
rect 1996 1470 2030 1486
rect 1996 1394 2030 1410
rect 2092 1470 2126 1486
rect 2092 1394 2126 1410
rect 2188 1470 2222 1486
rect 2188 1394 2222 1410
rect 2284 1470 2318 1486
rect 2284 1394 2318 1410
rect 2380 1470 2414 1486
rect 2380 1394 2414 1410
rect 2476 1470 2510 1486
rect 2476 1394 2510 1410
rect 2572 1470 2606 1486
rect 2572 1394 2606 1410
rect 2668 1470 2702 1486
rect 2668 1394 2702 1410
rect 2764 1470 2798 1486
rect 2764 1394 2798 1410
rect 2860 1470 2894 1486
rect 2860 1394 2894 1410
rect 2956 1470 2990 1486
rect 2956 1394 2990 1410
rect 3052 1470 3086 1486
rect 3052 1394 3086 1410
rect 3148 1470 3182 1486
rect 3148 1394 3182 1410
rect 3244 1470 3278 1486
rect 3244 1394 3278 1410
rect 3340 1470 3374 1486
rect 3340 1394 3374 1410
rect 3436 1470 3470 1486
rect 3436 1394 3470 1410
rect 3532 1470 3566 1486
rect 3532 1394 3566 1410
rect 3628 1470 3662 1486
rect 3628 1394 3662 1410
rect 3724 1470 3758 1486
rect 3724 1394 3758 1410
rect 3820 1470 3854 1486
rect 3820 1394 3854 1410
rect 3916 1470 3950 1486
rect 3916 1394 3950 1410
rect 4012 1470 4046 1486
rect 4012 1394 4046 1410
rect 4108 1470 4142 1486
rect 4108 1394 4142 1410
rect -1354 1366 -1262 1392
rect -1156 1324 1406 1360
rect 1548 1326 1564 1360
rect 1598 1326 1756 1360
rect 1790 1326 1948 1360
rect 1982 1326 2140 1360
rect 2174 1326 2332 1360
rect 2366 1326 2524 1360
rect 2558 1326 2716 1360
rect 2750 1326 2908 1360
rect 2942 1326 3100 1360
rect 3134 1326 3292 1360
rect 3326 1326 3484 1360
rect 3518 1326 3676 1360
rect 3710 1326 3868 1360
rect 3902 1326 4060 1360
rect 4094 1326 4110 1360
rect 1548 1324 4110 1326
<< viali >>
rect -1356 1978 -1312 2124
rect 1516 1872 1550 2100
rect 1612 1872 1646 2100
rect 1708 1872 1742 2100
rect 1804 1872 1838 2100
rect 1900 1872 1934 2100
rect 1996 1872 2030 2100
rect 2092 1872 2126 2100
rect 2188 1872 2222 2100
rect 2284 1872 2318 2100
rect 2380 1872 2414 2100
rect 2476 1872 2510 2100
rect 2572 1872 2606 2100
rect 2668 1872 2702 2100
rect 2764 1872 2798 2100
rect 2860 1872 2894 2100
rect 2956 1872 2990 2100
rect 3052 1872 3086 2100
rect 3148 1872 3182 2100
rect 3244 1872 3278 2100
rect 3340 1872 3374 2100
rect 3436 1872 3470 2100
rect 3532 1872 3566 2100
rect 3628 1872 3662 2100
rect 3724 1872 3758 2100
rect 3820 1872 3854 2100
rect 3916 1872 3950 2100
rect 4012 1872 4046 2100
rect 4108 1872 4142 2100
rect 1454 1564 1582 1666
rect -1336 1392 -1280 1456
rect 1516 1410 1550 1470
rect 1612 1410 1646 1470
rect 1708 1410 1742 1470
rect 1804 1410 1838 1470
rect 1900 1410 1934 1470
rect 1996 1410 2030 1470
rect 2092 1410 2126 1470
rect 2188 1410 2222 1470
rect 2284 1410 2318 1470
rect 2380 1410 2414 1470
rect 2476 1410 2510 1470
rect 2572 1410 2606 1470
rect 2668 1410 2702 1470
rect 2764 1410 2798 1470
rect 2860 1410 2894 1470
rect 2956 1410 2990 1470
rect 3052 1410 3086 1470
rect 3148 1410 3182 1470
rect 3244 1410 3278 1470
rect 3340 1410 3374 1470
rect 3436 1410 3470 1470
rect 3532 1410 3566 1470
rect 3628 1410 3662 1470
rect 3724 1410 3758 1470
rect 3820 1410 3854 1470
rect 3916 1410 3950 1470
rect 4012 1410 4046 1470
rect 4108 1410 4142 1470
<< metal1 >>
rect -1358 2260 -1118 2264
rect -1358 2230 1347 2260
rect -1358 2224 -1118 2230
rect -1356 2166 -1312 2224
rect -1378 2124 -1292 2166
rect -1378 1978 -1356 2124
rect -1312 1978 -1292 2124
rect -1188 2032 -1154 2224
rect -1104 2100 -1046 2112
rect -1378 1938 -1292 1978
rect -1048 1872 -1046 2100
rect -996 2028 -962 2230
rect -914 2100 -856 2112
rect -1104 1860 -1046 1872
rect -914 1872 -912 2100
rect -804 2038 -770 2230
rect -718 2100 -660 2112
rect -914 1860 -856 1872
rect -662 1872 -660 2100
rect -612 2036 -578 2230
rect -526 2100 -468 2112
rect -718 1860 -660 1872
rect -470 1872 -468 2100
rect -420 2040 -386 2230
rect -336 2100 -278 2112
rect -526 1860 -468 1872
rect -280 1872 -278 2100
rect -228 2034 -194 2230
rect -144 2100 -86 2112
rect -336 1860 -278 1872
rect -144 1872 -142 2100
rect -36 2032 -2 2230
rect 48 2100 106 2112
rect -144 1860 -86 1872
rect 48 1872 50 2100
rect 156 2032 190 2230
rect 240 2100 298 2112
rect 48 1860 106 1872
rect 296 1872 298 2100
rect 348 2028 382 2230
rect 432 2100 490 2114
rect 240 1860 298 1872
rect 488 1872 490 2100
rect 540 2024 574 2230
rect 626 2100 684 2114
rect 432 1862 490 1872
rect 682 1872 684 2100
rect 732 2038 766 2230
rect 816 2100 874 2112
rect 626 1862 684 1872
rect 816 1872 818 2100
rect 924 1990 958 2230
rect 1008 2100 1066 2112
rect 816 1860 874 1872
rect 1064 1872 1066 2100
rect 1116 1994 1150 2230
rect 1200 2100 1258 2112
rect 1008 1860 1066 1872
rect 1256 1872 1258 2100
rect 1317 1873 1347 2230
rect 1516 2230 4051 2260
rect 1516 2112 1550 2230
rect 1708 2112 1742 2230
rect 1900 2112 1934 2230
rect 2092 2112 2126 2230
rect 2284 2112 2318 2230
rect 2476 2112 2510 2230
rect 2668 2112 2702 2230
rect 2860 2112 2894 2230
rect 3052 2112 3086 2230
rect 1392 2100 1452 2112
rect 1200 1860 1258 1872
rect 1392 1872 1394 2100
rect 1450 1872 1452 2100
rect 1392 1862 1452 1872
rect 1510 2100 1556 2112
rect 1510 1872 1516 2100
rect 1550 1872 1556 2100
rect 1404 1682 1438 1862
rect 1510 1860 1556 1872
rect 1600 2100 1658 2112
rect 1656 1872 1658 2100
rect 1600 1860 1658 1872
rect 1702 2100 1748 2112
rect 1702 1872 1708 2100
rect 1742 1872 1748 2100
rect 1702 1860 1748 1872
rect 1790 2100 1848 2112
rect 1790 1872 1792 2100
rect 1790 1860 1848 1872
rect 1894 2100 1940 2112
rect 1894 1872 1900 2100
rect 1934 1872 1940 2100
rect 1894 1860 1940 1872
rect 1986 2100 2044 2112
rect 2042 1872 2044 2100
rect 1986 1860 2044 1872
rect 2086 2100 2132 2112
rect 2086 1872 2092 2100
rect 2126 1872 2132 2100
rect 2086 1860 2132 1872
rect 2178 2100 2236 2112
rect 2234 1872 2236 2100
rect 2178 1860 2236 1872
rect 2278 2100 2324 2112
rect 2278 1872 2284 2100
rect 2318 1872 2324 2100
rect 2278 1860 2324 1872
rect 2368 2100 2426 2112
rect 2424 1872 2426 2100
rect 2368 1860 2426 1872
rect 2470 2100 2516 2112
rect 2470 1872 2476 2100
rect 2510 1872 2516 2100
rect 2470 1860 2516 1872
rect 2560 2100 2618 2112
rect 2560 1872 2562 2100
rect 2560 1860 2618 1872
rect 2662 2100 2708 2112
rect 2662 1872 2668 2100
rect 2702 1872 2708 2100
rect 2662 1860 2708 1872
rect 2752 2100 2810 2112
rect 2752 1872 2754 2100
rect 2752 1860 2810 1872
rect 2854 2100 2900 2112
rect 2854 1872 2860 2100
rect 2894 1872 2900 2100
rect 2854 1860 2900 1872
rect 2944 2100 3002 2112
rect 3000 1872 3002 2100
rect 2944 1860 3002 1872
rect 3046 2100 3092 2112
rect 3046 1872 3052 2100
rect 3086 1872 3092 2100
rect 3046 1860 3092 1872
rect 3136 2100 3194 2114
rect 3244 2112 3278 2230
rect 3192 1872 3194 2100
rect 3136 1862 3194 1872
rect 3238 2100 3284 2112
rect 3238 1872 3244 2100
rect 3278 1872 3284 2100
rect 3142 1860 3188 1862
rect 3238 1860 3284 1872
rect 3330 2100 3388 2114
rect 3436 2112 3470 2230
rect 3628 2112 3662 2230
rect 3820 2112 3854 2230
rect 4021 2112 4051 2230
rect 3386 1872 3388 2100
rect 3330 1862 3388 1872
rect 3430 2100 3476 2112
rect 3430 1872 3436 2100
rect 3470 1872 3476 2100
rect 3334 1860 3380 1862
rect 3430 1860 3476 1872
rect 3520 2100 3578 2112
rect 3520 1872 3522 2100
rect 3520 1860 3578 1872
rect 3622 2100 3668 2112
rect 3622 1872 3628 2100
rect 3662 1872 3668 2100
rect 3622 1860 3668 1872
rect 3712 2100 3770 2112
rect 3768 1872 3770 2100
rect 3712 1860 3770 1872
rect 3814 2100 3860 2112
rect 3814 1872 3820 2100
rect 3854 1872 3860 2100
rect 3814 1860 3860 1872
rect 3904 2100 3962 2112
rect 3960 1872 3962 2100
rect 3904 1860 3962 1872
rect 4006 2100 4052 2112
rect 4006 1872 4012 2100
rect 4046 1872 4052 2100
rect 4006 1860 4052 1872
rect 4096 2100 4156 2112
rect 4096 1872 4098 2100
rect 4154 1872 4156 2100
rect 4096 1862 4156 1872
rect 4102 1860 4148 1862
rect 1404 1680 1476 1682
rect 1404 1666 1598 1680
rect 1404 1564 1454 1666
rect 1582 1564 1598 1666
rect 1404 1552 1598 1564
rect 1404 1484 1438 1552
rect 4108 1484 4142 1860
rect -1354 1456 -1262 1482
rect -1354 1392 -1336 1456
rect -1280 1392 -1262 1456
rect -1102 1470 -1044 1484
rect -1354 1366 -1262 1392
rect -1342 1304 -1270 1366
rect -1188 1305 -1154 1438
rect -1046 1410 -1044 1470
rect -910 1470 -852 1484
rect -1102 1398 -1044 1410
rect -996 1305 -962 1432
rect -854 1410 -852 1470
rect -720 1470 -662 1484
rect -910 1398 -852 1410
rect -804 1305 -770 1428
rect -664 1410 -662 1470
rect -528 1470 -470 1484
rect -720 1398 -662 1410
rect -612 1305 -578 1434
rect -472 1410 -470 1470
rect -338 1470 -280 1484
rect -528 1398 -470 1410
rect -420 1305 -386 1432
rect -338 1410 -336 1470
rect -144 1470 -86 1484
rect -338 1398 -280 1410
rect -228 1305 -194 1434
rect -88 1410 -86 1470
rect 48 1470 106 1484
rect -144 1398 -86 1410
rect -36 1305 -2 1432
rect 104 1410 106 1470
rect 242 1470 300 1484
rect 48 1398 106 1410
rect 156 1305 190 1430
rect 298 1410 300 1470
rect 434 1470 492 1484
rect 242 1398 300 1410
rect 348 1305 382 1436
rect 490 1410 492 1470
rect 624 1470 682 1484
rect 434 1398 492 1410
rect 540 1305 574 1434
rect 680 1410 682 1470
rect 818 1470 876 1484
rect 624 1398 682 1410
rect 732 1305 766 1432
rect 874 1410 876 1470
rect 1008 1470 1066 1484
rect 818 1398 876 1410
rect 924 1305 958 1434
rect 1064 1410 1066 1470
rect 1200 1470 1258 1484
rect 1008 1398 1066 1410
rect 1116 1305 1150 1434
rect 1256 1410 1258 1470
rect 1392 1470 1450 1484
rect 1200 1398 1258 1410
rect 1309 1305 1343 1423
rect 1448 1410 1450 1470
rect 1392 1398 1450 1410
rect 1510 1470 1556 1482
rect 1510 1410 1516 1470
rect 1550 1410 1556 1470
rect 1510 1398 1556 1410
rect 1602 1470 1660 1484
rect 1658 1410 1660 1470
rect 1602 1398 1660 1410
rect 1702 1470 1748 1482
rect 1702 1410 1708 1470
rect 1742 1410 1748 1470
rect 1702 1398 1748 1410
rect 1794 1470 1852 1484
rect 1850 1410 1852 1470
rect 1794 1398 1852 1410
rect 1894 1470 1940 1482
rect 1894 1410 1900 1470
rect 1934 1410 1940 1470
rect 1894 1398 1940 1410
rect 1984 1470 2042 1484
rect 2040 1410 2042 1470
rect 1984 1398 2042 1410
rect 2086 1470 2132 1482
rect 2086 1410 2092 1470
rect 2126 1410 2132 1470
rect 2086 1398 2132 1410
rect 2176 1470 2234 1484
rect 2232 1410 2234 1470
rect 2176 1398 2234 1410
rect 2278 1470 2324 1482
rect 2278 1410 2284 1470
rect 2318 1410 2324 1470
rect 2278 1398 2324 1410
rect 2366 1470 2424 1484
rect 2366 1410 2368 1470
rect 2366 1398 2424 1410
rect 2470 1470 2516 1482
rect 2470 1410 2476 1470
rect 2510 1410 2516 1470
rect 2470 1398 2516 1410
rect 2560 1470 2618 1484
rect 2616 1410 2618 1470
rect 2560 1398 2618 1410
rect 2662 1470 2708 1482
rect 2662 1410 2668 1470
rect 2702 1410 2708 1470
rect 2662 1398 2708 1410
rect 2752 1470 2810 1484
rect 2808 1410 2810 1470
rect 2752 1398 2810 1410
rect 2854 1470 2900 1482
rect 2854 1410 2860 1470
rect 2894 1410 2900 1470
rect 2854 1398 2900 1410
rect 2946 1470 3004 1484
rect 3002 1410 3004 1470
rect 2946 1398 3004 1410
rect 3046 1470 3092 1482
rect 3046 1410 3052 1470
rect 3086 1410 3092 1470
rect 3046 1398 3092 1410
rect 3138 1470 3196 1484
rect 3194 1410 3196 1470
rect 3138 1398 3196 1410
rect 3238 1470 3284 1482
rect 3238 1410 3244 1470
rect 3278 1410 3284 1470
rect 3238 1398 3284 1410
rect 3328 1470 3386 1484
rect 3384 1410 3386 1470
rect 3328 1398 3386 1410
rect 3430 1470 3476 1482
rect 3430 1410 3436 1470
rect 3470 1410 3476 1470
rect 3430 1398 3476 1410
rect 3522 1470 3580 1484
rect 3578 1410 3580 1470
rect 3522 1398 3580 1410
rect 3622 1470 3668 1482
rect 3622 1410 3628 1470
rect 3662 1410 3668 1470
rect 3622 1398 3668 1410
rect 3712 1470 3770 1484
rect 3768 1410 3770 1470
rect 3712 1398 3770 1410
rect 3814 1470 3860 1482
rect 3814 1410 3820 1470
rect 3854 1410 3860 1470
rect 3814 1398 3860 1410
rect 3904 1470 3962 1484
rect 3960 1410 3962 1470
rect 3904 1398 3962 1410
rect 4006 1470 4052 1482
rect 4006 1410 4012 1470
rect 4046 1410 4052 1470
rect 4006 1398 4052 1410
rect 4096 1470 4154 1484
rect 4152 1410 4154 1470
rect 4096 1398 4154 1410
rect -1188 1304 1343 1305
rect -1342 1274 1343 1304
rect -1188 1271 1343 1274
rect 1516 1305 1550 1398
rect 1708 1305 1742 1398
rect 1900 1305 1934 1398
rect 2092 1305 2126 1398
rect 2284 1305 2318 1398
rect 2476 1305 2510 1398
rect 2668 1305 2702 1398
rect 2860 1305 2894 1398
rect 3052 1305 3086 1398
rect 3244 1305 3278 1398
rect 3436 1305 3470 1398
rect 3628 1305 3662 1398
rect 3820 1305 3854 1398
rect 4013 1305 4047 1398
rect 1516 1271 4047 1305
<< via1 >>
rect -1104 1872 -1048 2100
rect -912 1872 -856 2100
rect -718 1872 -662 2100
rect -526 1872 -470 2100
rect -336 1872 -280 2100
rect -142 1872 -86 2100
rect 50 1872 106 2100
rect 240 1872 296 2100
rect 432 1872 488 2100
rect 626 1872 682 2100
rect 818 1872 874 2100
rect 1008 1872 1064 2100
rect 1200 1872 1256 2100
rect 1394 1872 1450 2100
rect 1600 1872 1612 2100
rect 1612 1872 1646 2100
rect 1646 1872 1656 2100
rect 1792 1872 1804 2100
rect 1804 1872 1838 2100
rect 1838 1872 1848 2100
rect 1986 1872 1996 2100
rect 1996 1872 2030 2100
rect 2030 1872 2042 2100
rect 2178 1872 2188 2100
rect 2188 1872 2222 2100
rect 2222 1872 2234 2100
rect 2368 1872 2380 2100
rect 2380 1872 2414 2100
rect 2414 1872 2424 2100
rect 2562 1872 2572 2100
rect 2572 1872 2606 2100
rect 2606 1872 2618 2100
rect 2754 1872 2764 2100
rect 2764 1872 2798 2100
rect 2798 1872 2810 2100
rect 2944 1872 2956 2100
rect 2956 1872 2990 2100
rect 2990 1872 3000 2100
rect 3136 1872 3148 2100
rect 3148 1872 3182 2100
rect 3182 1872 3192 2100
rect 3330 1872 3340 2100
rect 3340 1872 3374 2100
rect 3374 1872 3386 2100
rect 3522 1872 3532 2100
rect 3532 1872 3566 2100
rect 3566 1872 3578 2100
rect 3712 1872 3724 2100
rect 3724 1872 3758 2100
rect 3758 1872 3768 2100
rect 3904 1872 3916 2100
rect 3916 1872 3950 2100
rect 3950 1872 3960 2100
rect 4098 1872 4108 2100
rect 4108 1872 4142 2100
rect 4142 1872 4154 2100
rect -1102 1410 -1046 1470
rect -910 1410 -854 1470
rect -720 1410 -664 1470
rect -528 1410 -472 1470
rect -336 1410 -280 1470
rect -144 1410 -88 1470
rect 48 1410 104 1470
rect 242 1410 298 1470
rect 434 1410 490 1470
rect 624 1410 680 1470
rect 818 1410 874 1470
rect 1008 1410 1064 1470
rect 1200 1410 1256 1470
rect 1392 1410 1448 1470
rect 1602 1410 1612 1470
rect 1612 1410 1646 1470
rect 1646 1410 1658 1470
rect 1794 1410 1804 1470
rect 1804 1410 1838 1470
rect 1838 1410 1850 1470
rect 1984 1410 1996 1470
rect 1996 1410 2030 1470
rect 2030 1410 2040 1470
rect 2176 1410 2188 1470
rect 2188 1410 2222 1470
rect 2222 1410 2232 1470
rect 2368 1410 2380 1470
rect 2380 1410 2414 1470
rect 2414 1410 2424 1470
rect 2560 1410 2572 1470
rect 2572 1410 2606 1470
rect 2606 1410 2616 1470
rect 2752 1410 2764 1470
rect 2764 1410 2798 1470
rect 2798 1410 2808 1470
rect 2946 1410 2956 1470
rect 2956 1410 2990 1470
rect 2990 1410 3002 1470
rect 3138 1410 3148 1470
rect 3148 1410 3182 1470
rect 3182 1410 3194 1470
rect 3328 1410 3340 1470
rect 3340 1410 3374 1470
rect 3374 1410 3384 1470
rect 3522 1410 3532 1470
rect 3532 1410 3566 1470
rect 3566 1410 3578 1470
rect 3712 1410 3724 1470
rect 3724 1410 3758 1470
rect 3758 1410 3768 1470
rect 3904 1410 3916 1470
rect 3916 1410 3950 1470
rect 3950 1410 3960 1470
rect 4096 1410 4108 1470
rect 4108 1410 4142 1470
rect 4142 1410 4152 1470
<< metal2 >>
rect -1144 2100 1450 2112
rect -1144 1872 -1104 2100
rect -1048 1872 -912 2100
rect -856 1872 -718 2100
rect -662 1872 -526 2100
rect -470 1872 -336 2100
rect -280 1872 -142 2100
rect -86 1872 50 2100
rect 106 1872 240 2100
rect 296 1872 432 2100
rect 488 1872 626 2100
rect 682 1872 818 2100
rect 874 1872 1008 2100
rect 1064 1872 1200 2100
rect 1256 1872 1394 2100
rect -1144 1860 1450 1872
rect 1560 2100 4154 2112
rect 1560 1872 1600 2100
rect 1656 1872 1792 2100
rect 1848 1872 1986 2100
rect 2042 1872 2178 2100
rect 2234 1872 2368 2100
rect 2424 1872 2562 2100
rect 2618 1872 2754 2100
rect 2810 1872 2944 2100
rect 3000 1872 3136 2100
rect 3192 1872 3330 2100
rect 3386 1872 3522 2100
rect 3578 1872 3712 2100
rect 3768 1872 3904 2100
rect 3960 1872 4098 2100
rect 1560 1860 4154 1872
rect -1138 1470 1450 1484
rect -1138 1410 -1102 1470
rect -1046 1410 -910 1470
rect -854 1410 -720 1470
rect -664 1410 -528 1470
rect -472 1410 -336 1470
rect -280 1410 -144 1470
rect -88 1410 48 1470
rect 104 1410 242 1470
rect 298 1410 434 1470
rect 490 1410 624 1470
rect 680 1410 818 1470
rect 874 1410 1008 1470
rect 1064 1410 1200 1470
rect 1256 1410 1392 1470
rect 1448 1410 1450 1470
rect -1138 1398 1450 1410
rect 1566 1470 4154 1484
rect 1566 1410 1602 1470
rect 1658 1410 1794 1470
rect 1850 1410 1984 1470
rect 2040 1410 2176 1470
rect 2232 1410 2368 1470
rect 2424 1410 2560 1470
rect 2616 1410 2752 1470
rect 2808 1410 2946 1470
rect 3002 1410 3138 1470
rect 3194 1410 3328 1470
rect 3384 1410 3522 1470
rect 3578 1410 3712 1470
rect 3768 1410 3904 1470
rect 3960 1410 4096 1470
rect 4152 1410 4154 1470
rect 1566 1398 4154 1410
<< metal4 >>
rect -1330 2222 4170 2342
<< metal5 >>
rect -1320 776 4168 1314
use sky130_fd_pr__nfet_01v8_NJGLN5  sky130_fd_pr__nfet_01v8_NJGLN5_1
timestamp 1699103691
transform 1 0 125 0 1 1440
box -1325 -130 1325 130
use sky130_fd_pr__pfet_01v8_VR4B8J  sky130_fd_pr__pfet_01v8_VR4B8J_1
timestamp 1699103691
transform 1 0 125 0 1 1986
box -1361 -226 1361 226
<< end >>
