magic
tech sky130A
magscale 1 2
timestamp 1699103691
<< nmos >>
rect -687 -42 -657 42
rect -591 -42 -561 42
rect -495 -42 -465 42
rect -399 -42 -369 42
rect -303 -42 -273 42
rect -207 -42 -177 42
rect -111 -42 -81 42
rect -15 -42 15 42
rect 81 -42 111 42
rect 177 -42 207 42
rect 273 -42 303 42
rect 369 -42 399 42
rect 465 -42 495 42
rect 561 -42 591 42
rect 657 -42 687 42
<< ndiff >>
rect -749 30 -687 42
rect -749 -30 -737 30
rect -703 -30 -687 30
rect -749 -42 -687 -30
rect -657 30 -591 42
rect -657 -30 -641 30
rect -607 -30 -591 30
rect -657 -42 -591 -30
rect -561 30 -495 42
rect -561 -30 -545 30
rect -511 -30 -495 30
rect -561 -42 -495 -30
rect -465 30 -399 42
rect -465 -30 -449 30
rect -415 -30 -399 30
rect -465 -42 -399 -30
rect -369 30 -303 42
rect -369 -30 -353 30
rect -319 -30 -303 30
rect -369 -42 -303 -30
rect -273 30 -207 42
rect -273 -30 -257 30
rect -223 -30 -207 30
rect -273 -42 -207 -30
rect -177 30 -111 42
rect -177 -30 -161 30
rect -127 -30 -111 30
rect -177 -42 -111 -30
rect -81 30 -15 42
rect -81 -30 -65 30
rect -31 -30 -15 30
rect -81 -42 -15 -30
rect 15 30 81 42
rect 15 -30 31 30
rect 65 -30 81 30
rect 15 -42 81 -30
rect 111 30 177 42
rect 111 -30 127 30
rect 161 -30 177 30
rect 111 -42 177 -30
rect 207 30 273 42
rect 207 -30 223 30
rect 257 -30 273 30
rect 207 -42 273 -30
rect 303 30 369 42
rect 303 -30 319 30
rect 353 -30 369 30
rect 303 -42 369 -30
rect 399 30 465 42
rect 399 -30 415 30
rect 449 -30 465 30
rect 399 -42 465 -30
rect 495 30 561 42
rect 495 -30 511 30
rect 545 -30 561 30
rect 495 -42 561 -30
rect 591 30 657 42
rect 591 -30 607 30
rect 641 -30 657 30
rect 591 -42 657 -30
rect 687 30 749 42
rect 687 -30 703 30
rect 737 -30 749 30
rect 687 -42 749 -30
<< ndiffc >>
rect -737 -30 -703 30
rect -641 -30 -607 30
rect -545 -30 -511 30
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
rect 511 -30 545 30
rect 607 -30 641 30
rect 703 -30 737 30
<< poly >>
rect -609 114 -543 130
rect -609 80 -593 114
rect -559 80 -543 114
rect -687 42 -657 68
rect -609 64 -543 80
rect -417 114 -351 130
rect -417 80 -401 114
rect -367 80 -351 114
rect -591 42 -561 64
rect -495 42 -465 68
rect -417 64 -351 80
rect -225 114 -159 130
rect -225 80 -209 114
rect -175 80 -159 114
rect -399 42 -369 64
rect -303 42 -273 68
rect -225 64 -159 80
rect -33 114 33 130
rect -33 80 -17 114
rect 17 80 33 114
rect -207 42 -177 64
rect -111 42 -81 68
rect -33 64 33 80
rect 159 114 225 130
rect 159 80 175 114
rect 209 80 225 114
rect -15 42 15 64
rect 81 42 111 68
rect 159 64 225 80
rect 351 114 417 130
rect 351 80 367 114
rect 401 80 417 114
rect 177 42 207 64
rect 273 42 303 68
rect 351 64 417 80
rect 543 114 609 130
rect 543 80 559 114
rect 593 80 609 114
rect 369 42 399 64
rect 465 42 495 68
rect 543 64 609 80
rect 561 42 591 64
rect 657 42 687 68
rect -687 -64 -657 -42
rect -705 -80 -639 -64
rect -591 -68 -561 -42
rect -495 -64 -465 -42
rect -705 -114 -689 -80
rect -655 -114 -639 -80
rect -705 -130 -639 -114
rect -513 -80 -447 -64
rect -399 -68 -369 -42
rect -303 -64 -273 -42
rect -513 -114 -497 -80
rect -463 -114 -447 -80
rect -513 -130 -447 -114
rect -321 -80 -255 -64
rect -207 -68 -177 -42
rect -111 -64 -81 -42
rect -321 -114 -305 -80
rect -271 -114 -255 -80
rect -321 -130 -255 -114
rect -129 -80 -63 -64
rect -15 -68 15 -42
rect 81 -64 111 -42
rect -129 -114 -113 -80
rect -79 -114 -63 -80
rect -129 -130 -63 -114
rect 63 -80 129 -64
rect 177 -68 207 -42
rect 273 -64 303 -42
rect 63 -114 79 -80
rect 113 -114 129 -80
rect 63 -130 129 -114
rect 255 -80 321 -64
rect 369 -68 399 -42
rect 465 -64 495 -42
rect 255 -114 271 -80
rect 305 -114 321 -80
rect 255 -130 321 -114
rect 447 -80 513 -64
rect 561 -68 591 -42
rect 657 -64 687 -42
rect 447 -114 463 -80
rect 497 -114 513 -80
rect 447 -130 513 -114
rect 639 -80 705 -64
rect 639 -114 655 -80
rect 689 -114 705 -80
rect 639 -130 705 -114
<< polycont >>
rect -593 80 -559 114
rect -401 80 -367 114
rect -209 80 -175 114
rect -17 80 17 114
rect 175 80 209 114
rect 367 80 401 114
rect 559 80 593 114
rect -689 -114 -655 -80
rect -497 -114 -463 -80
rect -305 -114 -271 -80
rect -113 -114 -79 -80
rect 79 -114 113 -80
rect 271 -114 305 -80
rect 463 -114 497 -80
rect 655 -114 689 -80
<< locali >>
rect -609 80 -593 114
rect -559 80 -543 114
rect -417 80 -401 114
rect -367 80 -351 114
rect -225 80 -209 114
rect -175 80 -159 114
rect -33 80 -17 114
rect 17 80 33 114
rect 159 80 175 114
rect 209 80 225 114
rect 351 80 367 114
rect 401 80 417 114
rect 543 80 559 114
rect 593 80 609 114
rect -737 30 -703 46
rect -737 -46 -703 -30
rect -641 30 -607 46
rect -641 -46 -607 -30
rect -545 30 -511 46
rect -545 -46 -511 -30
rect -449 30 -415 46
rect -449 -46 -415 -30
rect -353 30 -319 46
rect -353 -46 -319 -30
rect -257 30 -223 46
rect -257 -46 -223 -30
rect -161 30 -127 46
rect -161 -46 -127 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 127 30 161 46
rect 127 -46 161 -30
rect 223 30 257 46
rect 223 -46 257 -30
rect 319 30 353 46
rect 319 -46 353 -30
rect 415 30 449 46
rect 415 -46 449 -30
rect 511 30 545 46
rect 511 -46 545 -30
rect 607 30 641 46
rect 607 -46 641 -30
rect 703 30 737 46
rect 703 -46 737 -30
rect -705 -114 -689 -80
rect -655 -114 -639 -80
rect -513 -114 -497 -80
rect -463 -114 -447 -80
rect -321 -114 -305 -80
rect -271 -114 -255 -80
rect -129 -114 -113 -80
rect -79 -114 -63 -80
rect 63 -114 79 -80
rect 113 -114 129 -80
rect 255 -114 271 -80
rect 305 -114 321 -80
rect 447 -114 463 -80
rect 497 -114 513 -80
rect 639 -114 655 -80
rect 689 -114 705 -80
<< viali >>
rect -737 -30 -703 30
rect -641 -30 -607 30
rect -545 -30 -511 30
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
rect 511 -30 545 30
rect 607 -30 641 30
rect 703 -30 737 30
<< metal1 >>
rect -743 30 -697 42
rect -743 -30 -737 30
rect -703 -30 -697 30
rect -743 -42 -697 -30
rect -647 30 -601 42
rect -647 -30 -641 30
rect -607 -30 -601 30
rect -647 -42 -601 -30
rect -551 30 -505 42
rect -551 -30 -545 30
rect -511 -30 -505 30
rect -551 -42 -505 -30
rect -455 30 -409 42
rect -455 -30 -449 30
rect -415 -30 -409 30
rect -455 -42 -409 -30
rect -359 30 -313 42
rect -359 -30 -353 30
rect -319 -30 -313 30
rect -359 -42 -313 -30
rect -263 30 -217 42
rect -263 -30 -257 30
rect -223 -30 -217 30
rect -263 -42 -217 -30
rect -167 30 -121 42
rect -167 -30 -161 30
rect -127 -30 -121 30
rect -167 -42 -121 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 121 30 167 42
rect 121 -30 127 30
rect 161 -30 167 30
rect 121 -42 167 -30
rect 217 30 263 42
rect 217 -30 223 30
rect 257 -30 263 30
rect 217 -42 263 -30
rect 313 30 359 42
rect 313 -30 319 30
rect 353 -30 359 30
rect 313 -42 359 -30
rect 409 30 455 42
rect 409 -30 415 30
rect 449 -30 455 30
rect 409 -42 455 -30
rect 505 30 551 42
rect 505 -30 511 30
rect 545 -30 551 30
rect 505 -42 551 -30
rect 601 30 647 42
rect 601 -30 607 30
rect 641 -30 647 30
rect 601 -42 647 -30
rect 697 30 743 42
rect 697 -30 703 30
rect 737 -30 743 30
rect 697 -42 743 -30
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 15 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
