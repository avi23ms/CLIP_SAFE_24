* SPICE3 file created from capacitors.ext - technology: sky130A

X0 capacitor_7_0/buffer_and_gate_0/clk_out m3_n90_n15462# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1 capacitor_7_1/buffer_and_gate_0/clk_out m3_n90_n15462# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X2 capacitor_7_2/buffer_and_gate_0/clk_out m3_n90_n15462# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X3 capacitor_7_3/buffer_and_gate_0/clk_out m3_n90_n15462# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X4 capacitor_7_4/buffer_and_gate_0/clk_out m3_n90_n15462# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X5 capacitor_7_5/buffer_and_gate_0/clk_out m3_n90_n15462# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X6 capacitor_7_6/buffer_and_gate_0/clk_out m3_n90_n15462# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X7 capacitor_7_7/buffer_and_gate_0/clk_out m3_n90_n15462# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
C0 capacitor_7_3/buffer_and_gate_0/vdd capacitor_7_3/buffer_and_gate_0/m1_5444_838# 8.43f
C1 capacitor_7_2/buffer_and_gate_0/m1_5444_838# capacitor_7_2/buffer_and_gate_0/buffer_0/a_1436_1552# 2.15f
C2 capacitor_7_1/buffer_and_gate_0/vdd VSUBS 10.9f
C3 capacitor_7_5/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_5/buffer_and_gate_0/m1_5444_838# 2.15f
C4 capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 3.96f
C5 capacitor_7_6/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_6/buffer_and_gate_0/clk 2.22f
C6 capacitor_7_4/buffer_and_gate_0/and_gate_0/a_n78_396# capacitor_7_4/buffer_and_gate_0/vdd 3.45f
C7 capacitor_7_2/buffer_and_gate_0/m1_5444_838# VSUBS 4.04f
C8 capacitor_7_3/buffer_and_gate_0/vdd VSUBS 10.9f
C9 capacitor_7_3/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_3/buffer_and_gate_0/clk 2.22f
C10 capacitor_7_5/buffer_and_gate_0/m1_5444_838# VSUBS 4.04f
C11 capacitor_7_6/buffer_and_gate_0/clk capacitor_7_6/buffer_and_gate_0/vdd 4.6f
C12 capacitor_7_6/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.01f
C13 VSUBS capacitor_7_4/buffer_and_gate_0/vdd 11f
C14 capacitor_7_2/buffer_and_gate_0/vdd capacitor_7_2/buffer_and_gate_0/buffer_0/a_1436_1552# 12.9f
C15 capacitor_7_7/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_7/buffer_and_gate_0/clk 2.22f
C16 capacitor_7_0/buffer_and_gate_0/m1_5444_838# capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.15f
C17 capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 5.87f
C18 capacitor_7_2/buffer_and_gate_0/vdd capacitor_7_2/buffer_and_gate_0/and_gate_0/a_n78_396# 3.45f
C19 capacitor_7_0/buffer_and_gate_0/m1_5444_838# capacitor_7_0/buffer_and_gate_0/vdd 8.43f
C20 capacitor_7_6/buffer_and_gate_0/vdd VSUBS 10.4f
C21 capacitor_7_2/buffer_and_gate_0/vdd capacitor_7_2/buffer_and_gate_0/clk 4.6f
C22 capacitor_7_2/buffer_and_gate_0/vdd VSUBS 10.9f
C23 capacitor_7_1/buffer_and_gate_0/vdd capacitor_7_1/buffer_and_gate_0/buffer_0/a_1436_1552# 12.9f
C24 capacitor_7_1/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.01f
C25 capacitor_7_3/buffer_and_gate_0/vdd capacitor_7_3/buffer_and_gate_0/and_gate_0/a_n78_396# 3.45f
C26 capacitor_7_2/buffer_and_gate_0/vdd capacitor_7_2/buffer_and_gate_0/m1_5444_838# 8.43f
C27 capacitor_7_6/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_6/buffer_and_gate_0/vdd 12.9f
C28 capacitor_7_7/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_7/buffer_and_gate_0/vdd 12.9f
C29 capacitor_7_7/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_7/buffer_and_gate_0/m1_5444_838# 2.15f
C30 capacitor_7_0/buffer_and_gate_0/vdd capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 12.9f
C31 capacitor_7_4/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.01f
C32 capacitor_7_4/buffer_and_gate_0/m1_5444_838# VSUBS 4.04f
C33 capacitor_7_7/buffer_and_gate_0/vdd VSUBS 10.9f
C34 capacitor_7_7/buffer_and_gate_0/m1_5444_838# VSUBS 4.04f
C35 capacitor_7_5/buffer_and_gate_0/clk capacitor_7_5/buffer_and_gate_0/vdd 4.6f
C36 capacitor_7_5/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_5/buffer_and_gate_0/vdd 12.9f
C37 capacitor_7_1/buffer_and_gate_0/vdd capacitor_7_1/buffer_and_gate_0/clk 4.6f
C38 capacitor_7_3/buffer_and_gate_0/m1_5444_838# capacitor_7_3/buffer_and_gate_0/buffer_0/a_1436_1552# 2.15f
C39 capacitor_7_3/buffer_and_gate_0/vdd capacitor_7_3/buffer_and_gate_0/clk 4.6f
C40 capacitor_7_1/buffer_and_gate_0/vdd capacitor_7_1/buffer_and_gate_0/m1_5444_838# 8.43f
C41 capacitor_7_5/buffer_and_gate_0/and_gate_0/a_n78_396# capacitor_7_5/buffer_and_gate_0/vdd 3.45f
C42 capacitor_7_4/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_4/buffer_and_gate_0/vdd 12.9f
C43 capacitor_7_1/buffer_and_gate_0/m1_5444_838# VSUBS 4.04f
C44 capacitor_7_4/buffer_and_gate_0/m1_5444_838# capacitor_7_4/buffer_and_gate_0/vdd 8.43f
C45 capacitor_7_5/buffer_and_gate_0/vdd VSUBS 10.9f
C46 capacitor_7_6/buffer_and_gate_0/and_gate_0/a_n78_396# capacitor_7_6/buffer_and_gate_0/vdd 3.45f
C47 capacitor_7_3/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.01f
C48 capacitor_7_4/buffer_and_gate_0/clk capacitor_7_4/buffer_and_gate_0/vdd 4.6f
C49 capacitor_7_7/buffer_and_gate_0/vdd capacitor_7_7/buffer_and_gate_0/clk 4.6f
C50 capacitor_7_5/buffer_and_gate_0/m1_5444_838# capacitor_7_5/buffer_and_gate_0/vdd 8.43f
C51 capacitor_7_6/buffer_and_gate_0/m1_5444_838# VSUBS 4.04f
C52 capacitor_7_3/buffer_and_gate_0/vdd capacitor_7_3/buffer_and_gate_0/buffer_0/a_1436_1552# 12.9f
C53 capacitor_7_1/buffer_and_gate_0/clk capacitor_7_1/buffer_and_gate_0/buffer_0/a_1436_1552# 2.22f
C54 capacitor_7_5/buffer_and_gate_0/clk capacitor_7_5/buffer_and_gate_0/buffer_0/a_1436_1552# 2.22f
C55 capacitor_7_6/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_6/buffer_and_gate_0/m1_5444_838# 2.15f
C56 capacitor_7_1/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_1/buffer_and_gate_0/m1_5444_838# 2.15f
C57 capacitor_7_4/buffer_and_gate_0/m1_5444_838# capacitor_7_4/buffer_and_gate_0/buffer_0/a_1436_1552# 2.15f
C58 capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# capacitor_7_0/buffer_and_gate_0/clk 2.22f
C59 capacitor_7_1/buffer_and_gate_0/vdd capacitor_7_1/buffer_and_gate_0/and_gate_0/a_n78_396# 3.45f
C60 capacitor_7_0/buffer_and_gate_0/vdd capacitor_7_0/buffer_and_gate_0/clk 4.6f
C61 capacitor_7_7/buffer_and_gate_0/vdd capacitor_7_7/buffer_and_gate_0/and_gate_0/a_n78_396# 3.45f
C62 capacitor_7_7/buffer_and_gate_0/vdd capacitor_7_7/buffer_and_gate_0/m1_5444_838# 8.43f
C63 capacitor_7_6/buffer_and_gate_0/vdd capacitor_7_6/buffer_and_gate_0/m1_5444_838# 8.43f
C64 capacitor_7_3/buffer_and_gate_0/m1_5444_838# VSUBS 4.04f
C65 capacitor_7_0/buffer_and_gate_0/vdd capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.45f
C66 capacitor_7_4/buffer_and_gate_0/clk capacitor_7_4/buffer_and_gate_0/buffer_0/a_1436_1552# 2.22f
C67 capacitor_7_2/buffer_and_gate_0/clk capacitor_7_2/buffer_and_gate_0/buffer_0/a_1436_1552# 2.22f
C68 capacitor_7_5/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.01f
C69 capacitor_7_7/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.01f
C70 capacitor_7_2/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.01f
Xcapacitor_7_0/buffer_and_gate_0 capacitor_7_0/buffer_and_gate_0/vdd VSUBS capacitor_7_0/buffer_and_gate_0/in
+ capacitor_7_0/buffer_and_gate_0/clk capacitor_7_0/buffer_and_gate_0/clk_out buffer_and_gate
Xcapacitor_7_1/buffer_and_gate_0 capacitor_7_1/buffer_and_gate_0/vdd VSUBS capacitor_7_1/buffer_and_gate_0/in
+ capacitor_7_1/buffer_and_gate_0/clk capacitor_7_1/buffer_and_gate_0/clk_out buffer_and_gate
Xcapacitor_7_2/buffer_and_gate_0 capacitor_7_2/buffer_and_gate_0/vdd VSUBS capacitor_7_2/buffer_and_gate_0/in
+ capacitor_7_2/buffer_and_gate_0/clk capacitor_7_2/buffer_and_gate_0/clk_out buffer_and_gate
Xcapacitor_7_3/buffer_and_gate_0 capacitor_7_3/buffer_and_gate_0/vdd VSUBS capacitor_7_3/buffer_and_gate_0/in
+ capacitor_7_3/buffer_and_gate_0/clk capacitor_7_3/buffer_and_gate_0/clk_out buffer_and_gate
Xcapacitor_7_4/buffer_and_gate_0 capacitor_7_4/buffer_and_gate_0/vdd VSUBS capacitor_7_4/buffer_and_gate_0/in
+ capacitor_7_4/buffer_and_gate_0/clk capacitor_7_4/buffer_and_gate_0/clk_out buffer_and_gate
Xcapacitor_7_5/buffer_and_gate_0 capacitor_7_5/buffer_and_gate_0/vdd VSUBS capacitor_7_5/buffer_and_gate_0/in
+ capacitor_7_5/buffer_and_gate_0/clk capacitor_7_5/buffer_and_gate_0/clk_out buffer_and_gate
Xcapacitor_7_6/buffer_and_gate_0 capacitor_7_6/buffer_and_gate_0/vdd VSUBS capacitor_7_6/buffer_and_gate_0/in
+ capacitor_7_6/buffer_and_gate_0/clk capacitor_7_6/buffer_and_gate_0/clk_out buffer_and_gate
Xcapacitor_7_7/buffer_and_gate_0 capacitor_7_7/buffer_and_gate_0/vdd VSUBS capacitor_7_7/buffer_and_gate_0/in
+ capacitor_7_7/buffer_and_gate_0/clk capacitor_7_7/buffer_and_gate_0/clk_out buffer_and_gate
C71 m3_n90_n15462# 0 16.3f **FLOATING
C72 capacitor_7_7/buffer_and_gate_0/in 0 3.04f
C73 capacitor_7_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.31f
C74 capacitor_7_7/buffer_and_gate_0/clk 0 7.7f
C75 capacitor_7_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C76 capacitor_7_7/buffer_and_gate_0/vdd 0 17.6f
C77 VSUBS 0 57.4f
C78 capacitor_7_6/buffer_and_gate_0/in 0 3.04f
C79 capacitor_7_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.31f
C80 capacitor_7_6/buffer_and_gate_0/clk 0 7.7f
C81 capacitor_7_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C82 capacitor_7_6/buffer_and_gate_0/vdd 0 17.6f
C83 capacitor_7_5/buffer_and_gate_0/in 0 3.04f
C84 capacitor_7_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.31f
C85 capacitor_7_5/buffer_and_gate_0/clk 0 7.7f
C86 capacitor_7_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C87 capacitor_7_5/buffer_and_gate_0/vdd 0 17.6f
C88 capacitor_7_4/buffer_and_gate_0/in 0 3.04f
C89 capacitor_7_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.31f
C90 capacitor_7_4/buffer_and_gate_0/clk 0 7.7f
C91 capacitor_7_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C92 capacitor_7_4/buffer_and_gate_0/vdd 0 17.6f
C93 capacitor_7_3/buffer_and_gate_0/in 0 3.04f
C94 capacitor_7_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.31f
C95 capacitor_7_3/buffer_and_gate_0/clk 0 7.7f
C96 capacitor_7_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C97 capacitor_7_3/buffer_and_gate_0/vdd 0 17.6f
C98 capacitor_7_2/buffer_and_gate_0/in 0 3.04f
C99 capacitor_7_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.31f
C100 capacitor_7_2/buffer_and_gate_0/clk 0 7.7f
C101 capacitor_7_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C102 capacitor_7_2/buffer_and_gate_0/vdd 0 17.6f
C103 capacitor_7_1/buffer_and_gate_0/in 0 3.04f
C104 capacitor_7_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.31f
C105 capacitor_7_1/buffer_and_gate_0/clk 0 7.7f
C106 capacitor_7_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C107 capacitor_7_1/buffer_and_gate_0/vdd 0 17.6f
C108 capacitor_7_0/buffer_and_gate_0/in 0 3.04f
C109 capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.31f
C110 capacitor_7_0/buffer_and_gate_0/clk 0 7.7f
C111 capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C112 capacitor_7_0/buffer_and_gate_0/vdd 0 17.6f
