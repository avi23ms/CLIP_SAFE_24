magic
tech sky130A
magscale 1 2
timestamp 1698488976
<< dnwell >>
rect 118 -1078 1558 -38
<< nwell >>
rect 12 -66 1674 102
rect 12 -78 1672 -66
rect 12 -1012 272 -78
rect 1424 -1012 1672 -78
rect 12 -1196 1672 -1012
rect 12 -1198 260 -1196
rect 1424 -1200 1672 -1196
<< nsubdiff >>
rect 88 -682 202 -656
rect 88 -966 112 -682
rect 180 -966 202 -682
rect 1488 -678 1602 -650
rect 88 -990 202 -966
rect 1488 -960 1510 -678
rect 1576 -960 1602 -678
rect 1488 -984 1602 -960
<< nsubdiffcont >>
rect 112 -966 180 -682
rect 1510 -960 1576 -678
<< poly >>
rect 410 -824 610 -764
rect 1028 -822 1228 -770
rect 1020 -824 1228 -822
rect 410 -840 630 -824
rect 410 -876 442 -840
rect 608 -876 630 -840
rect 410 -892 630 -876
rect 1008 -840 1228 -824
rect 1008 -874 1026 -840
rect 1186 -874 1228 -840
rect 1008 -892 1228 -874
<< polycont >>
rect 442 -876 608 -840
rect 1026 -874 1186 -840
<< locali >>
rect 88 -682 202 -656
rect 88 -966 112 -682
rect 180 -966 202 -682
rect 1488 -678 1602 -650
rect 1020 -824 1228 -822
rect 410 -840 630 -824
rect 410 -876 442 -840
rect 608 -876 630 -840
rect 410 -892 630 -876
rect 1008 -840 1228 -824
rect 1008 -874 1026 -840
rect 1186 -874 1228 -840
rect 1008 -892 1228 -874
rect 88 -990 202 -966
rect 1488 -960 1510 -678
rect 1576 -960 1602 -678
rect 1488 -984 1602 -960
<< viali >>
rect 112 -966 180 -682
rect 442 -876 608 -840
rect 1026 -874 1186 -840
rect 1510 -960 1576 -678
<< metal1 >>
rect 88 -682 202 -656
rect 88 -966 112 -682
rect 180 -936 202 -682
rect 1488 -678 1602 -650
rect 362 -766 400 -702
rect 364 -935 398 -766
rect 622 -824 656 -742
rect 982 -824 1016 -742
rect 1239 -766 1277 -711
rect 426 -840 1208 -824
rect 426 -876 442 -840
rect 608 -874 1026 -840
rect 1186 -874 1208 -840
rect 608 -876 1208 -874
rect 426 -892 1208 -876
rect 1239 -884 1273 -766
rect 1239 -934 1272 -884
rect 1488 -934 1510 -678
rect 1238 -935 1510 -934
rect 364 -936 1510 -935
rect 180 -960 1510 -936
rect 1576 -960 1602 -678
rect 180 -966 1602 -960
rect 88 -969 1602 -966
rect 88 -972 440 -969
rect 1238 -970 1602 -969
rect 88 -990 202 -972
rect 1488 -984 1602 -970
use sky130_fd_pr__nfet_01v8_EFUU27  sky130_fd_pr__nfet_01v8_EFUU27_0
timestamp 1698341146
transform 1 0 1128 0 1 -462
box -158 -326 158 326
use sky130_fd_pr__nfet_01v8_EFUU27  sky130_fd_pr__nfet_01v8_EFUU27_1
timestamp 1698341146
transform 1 0 510 0 1 -464
box -158 -326 158 326
<< end >>
