magic
tech sky130A
magscale 1 2
timestamp 1727007906
<< psubdiff >>
rect 384 2722 910 2806
rect 384 2554 446 2722
rect 814 2554 910 2722
rect 384 2486 910 2554
<< psubdiffcont >>
rect 446 2554 814 2722
<< poly >>
rect 696 3302 834 3316
rect 696 3244 722 3302
rect 806 3244 834 3302
rect 696 3230 834 3244
rect 712 3162 812 3230
<< polycont >>
rect 722 3244 806 3302
<< locali >>
rect 696 3302 834 3316
rect 696 3244 722 3302
rect 806 3244 834 3302
rect 696 3230 834 3244
rect 384 2722 910 2806
rect 384 2554 446 2722
rect 814 2554 910 2722
rect 384 2486 910 2554
<< viali >>
rect 722 3244 806 3302
rect 446 2554 814 2722
<< metal1 >>
rect 2582 4618 2746 4636
rect 2582 4546 2608 4618
rect 2720 4546 2746 4618
rect 2582 4524 2746 4546
rect 592 3478 636 3484
rect 572 3454 636 3478
rect 572 3156 616 3454
rect 697 3316 3060 3326
rect 696 3302 3060 3316
rect 696 3244 722 3302
rect 806 3276 3060 3302
rect 806 3244 834 3276
rect 696 3230 834 3244
rect 572 3118 698 3156
rect 572 2806 616 3118
rect 1015 3111 1065 3276
rect 2508 3228 2826 3240
rect 2508 3222 2848 3228
rect 2508 3164 2552 3222
rect 2816 3168 2848 3222
rect 2816 3164 2826 3168
rect 2508 3150 2826 3164
rect 827 3061 1065 3111
rect 384 2722 910 2806
rect 384 2554 446 2722
rect 814 2554 910 2722
rect 384 2486 910 2554
<< via1 >>
rect 2608 4546 2720 4618
rect 2552 3164 2816 3222
<< metal2 >>
rect 2582 4618 2746 4636
rect 2582 4546 2608 4618
rect 2720 4546 2746 4618
rect 2582 4524 2746 4546
rect 2508 3228 2826 3240
rect 2508 3222 2848 3228
rect 2508 3164 2552 3222
rect 2816 3168 2848 3222
rect 2816 3164 2826 3168
rect 2508 3150 2826 3164
<< via2 >>
rect 2608 4546 2720 4618
rect 2552 3164 2816 3222
<< metal3 >>
rect 2558 4618 2784 4640
rect 2558 4546 2608 4618
rect 2720 4546 2784 4618
rect 2558 4516 2784 4546
rect 2622 3240 2720 4516
rect 2508 3228 2826 3240
rect 2508 3222 2848 3228
rect 2508 3164 2552 3222
rect 2816 3168 2848 3222
rect 2816 3164 2826 3168
rect 2508 3150 2826 3164
use integrator_full_new_compact  integrator_full_new_compact_0
timestamp 1698861754
transform 1 0 394 0 1 3504
box -386 -3496 4003 1133
use sky130_fd_pr__nfet_01v8_LYF9NA  sky130_fd_pr__nfet_01v8_LYF9NA_0
timestamp 1726930802
transform 1 0 762 0 1 3046
box -108 -126 108 126
<< labels >>
rlabel metal1 1124 3300 1124 3300 1 vbias_integrator
<< end >>
