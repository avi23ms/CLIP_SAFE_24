magic
tech sky130A
magscale 1 2
timestamp 1698474034
<< metal1 >>
rect 7467 3015 7501 4220
rect 15136 3070 15481 3104
rect 7467 2981 8039 3015
rect 7467 863 7501 2981
rect 16798 962 18110 1006
rect 16798 954 16824 962
rect 14883 920 16824 954
rect 7467 829 7821 863
rect 16798 830 16824 920
rect 17226 830 18110 962
rect 7467 116 7501 829
rect 16798 798 18110 830
rect 7297 82 7501 116
rect 7332 -60 7480 -24
rect 7444 -1374 7480 -60
rect 16796 -1238 17996 -1206
rect 16796 -1298 16872 -1238
rect 14864 -1332 16872 -1298
rect 16796 -1368 16872 -1332
rect 17136 -1368 17996 -1238
rect 7444 -1410 7888 -1374
rect 7444 -3492 7480 -1410
rect 16796 -1416 17996 -1368
rect 14897 -3416 15325 -3382
rect 7444 -3528 7782 -3492
rect 7444 -4326 7480 -3528
<< via1 >>
rect 16824 830 17226 962
rect 16872 -1368 17136 -1238
<< metal2 >>
rect 7410 3120 7988 3160
rect 7410 -946 7450 3120
rect 7414 -1666 7450 -946
rect 7536 958 7724 998
rect 7536 -1254 7576 958
rect 7536 -1294 7920 -1254
rect 7410 -3338 7450 -1666
rect 7410 -3378 7734 -3338
rect 15628 -4326 15668 4220
rect 16798 962 17306 1004
rect 16798 830 16824 962
rect 17226 830 17306 962
rect 16798 798 17306 830
rect 16796 -1238 17198 -1202
rect 16796 -1368 16872 -1238
rect 17136 -1368 17198 -1238
rect 16796 -1416 17198 -1368
<< via2 >>
rect 16824 830 17226 962
rect 16872 -1368 17136 -1238
<< metal3 >>
rect 16798 962 17306 1004
rect 16798 830 16824 962
rect 17226 830 17306 962
rect 16798 798 17306 830
rect 18930 592 19396 806
rect 1014 68 1244 160
rect 16796 -1238 17198 -1202
rect 16796 -1368 16872 -1238
rect 17136 -1368 17198 -1238
rect 16796 -1416 17198 -1368
rect 18576 -1396 19540 -1196
<< via3 >>
rect 16824 830 17226 962
rect 16872 -1368 17136 -1238
<< metal4 >>
rect 15620 3976 15804 4220
rect 14734 3792 15804 3976
rect 7208 1952 15518 1996
rect 15620 1952 15804 3792
rect 7208 1812 15804 1952
rect 7208 954 7392 1812
rect 15334 1768 15804 1812
rect 15334 -396 15518 1768
rect 14304 -580 15518 -396
rect 15620 -2446 15804 1768
rect 16798 962 18110 1006
rect 16798 830 16824 962
rect 17226 830 18110 962
rect 16798 798 18110 830
rect 16796 -1238 17996 -1206
rect 16796 -1368 16872 -1238
rect 17136 -1368 17996 -1238
rect 16796 -1416 17996 -1368
rect 14538 -2630 15804 -2446
rect 15566 -4326 15750 -2630
<< metal5 >>
rect 15773 3070 16343 4220
rect 15784 2728 16343 3070
rect 14702 2671 16343 2728
rect 14697 2101 16343 2671
rect 15773 580 16343 2101
rect 15019 452 16343 580
rect 14428 76 16343 452
rect 15019 10 16343 76
rect 6736 -1034 6950 -1030
rect 6966 -1034 7350 -996
rect 6736 -1036 7350 -1034
rect 6720 -1556 7350 -1036
rect 6720 -1666 7362 -1556
rect 6720 -1828 7970 -1666
rect 15400 -1672 16343 10
rect 14992 -1828 16343 -1672
rect 6720 -2204 16343 -1828
rect 6966 -2212 7970 -2204
rect 14992 -2242 16343 -2204
rect 15444 -2244 16343 -2242
rect 15773 -3735 16343 -2244
rect 14683 -4305 16343 -3735
rect 15773 -4326 16343 -4305
use buffer_and_gate  buffer_and_gate_0
timestamp 1698472463
transform 1 0 7758 0 1 40
box -116 -30 7470 2020
use buffer_and_gate  buffer_and_gate_1
timestamp 1698472463
transform 1 0 7736 0 1 -2212
box -116 -30 7470 2020
use buffer_and_gate  buffer_and_gate_2
timestamp 1698472463
transform 1 0 8008 0 1 2190
box -116 -30 7470 2020
use buffer_and_gate  buffer_and_gate_3
timestamp 1698472463
transform 1 0 7774 0 1 -4296
box -116 -30 7470 2020
use clock  clock_0
timestamp 1698410772
transform 1 0 1368 0 1 216
box -410 -1832 6030 1274
use sky130_fd_pr__cap_mim_m3_1_VEQCNX  sky130_fd_pr__cap_mim_m3_1_VEQCNX_0
timestamp 0
transform 1 0 18280 0 1 742
box -886 -740 886 740
use sky130_fd_pr__cap_mim_m3_1_VEQCNX  sky130_fd_pr__cap_mim_m3_1_VEQCNX_1
timestamp 0
transform 1 0 18282 0 1 -1458
box -886 -740 886 740
<< labels >>
rlabel metal3 1052 106 1052 106 1 clk_in
port 1 n
rlabel space 1784 1132 1784 1132 1 vdd
port 2 n
rlabel metal4 7326 1688 7326 1688 1 vdd
port 3 n
rlabel metal5 7326 -2058 7326 -2058 1 gnd
port 4 n
rlabel metal1 7490 584 7490 584 1 clk
port 5 n
rlabel metal1 7462 -264 7462 -264 1 clkb
port 6 n
rlabel metal2 7600 974 7600 974 1 in1
port 7 n
rlabel metal1 15122 -1318 15122 -1318 1 clkb_out
port 8 n
rlabel metal1 15054 932 15054 932 1 clk_out
port 9 n
rlabel metal2 7602 -3376 7602 -3376 1 in2
port 11 n
rlabel metal1 15404 3082 15404 3082 1 clk2
port 13 n
rlabel metal1 15248 -3398 15248 -3398 1 clkb2
port 14 n
rlabel metal3 19308 714 19308 714 1 cap1
port 23 n
rlabel metal3 19448 -1300 19448 -1300 1 cap2
port 24 n
<< end >>
