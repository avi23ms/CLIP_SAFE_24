magic
tech sky130A
magscale 1 2
timestamp 1698861754
<< locali >>
rect 3212 -64 3618 -50
rect 3212 -120 3700 -64
<< metal1 >>
rect 192 1061 392 1102
rect 2896 1022 3616 1116
rect 1946 216 1956 304
rect 2032 216 2042 304
rect 514 118 524 176
rect 628 118 638 176
rect 888 164 1050 178
rect 888 112 918 164
rect 1020 112 1050 164
rect 3488 148 3504 166
rect 888 90 1050 112
rect 3364 -42 3618 10
rect 2968 -220 3154 -186
rect 2968 -268 3156 -220
rect 2968 -304 3604 -268
rect 1702 -598 1712 -500
rect 1778 -598 1788 -500
<< via1 >>
rect 1956 216 2032 304
rect 524 118 628 176
rect 918 112 1020 164
rect 1712 -598 1778 -500
<< metal2 >>
rect 1966 314 2002 346
rect 1956 312 2032 314
rect 1948 304 2040 312
rect 1948 216 1956 304
rect 2032 216 2040 304
rect 1948 200 2040 216
rect 540 186 606 188
rect 524 176 628 186
rect 932 174 978 178
rect 918 172 1020 174
rect 524 108 628 118
rect 910 164 1046 172
rect 910 112 918 164
rect 1020 112 1046 164
rect 540 -1269 606 108
rect 910 96 1046 112
rect 932 -119 978 96
rect 932 -165 1765 -119
rect 1719 -480 1765 -165
rect 1966 -276 2002 200
rect 1828 -278 2002 -276
rect 1826 -314 2002 -278
rect 1710 -500 1782 -480
rect 1710 -592 1712 -500
rect 1778 -592 1782 -500
rect 1826 -546 1864 -314
rect 1712 -608 1778 -598
rect 1826 -696 1862 -546
use cmfb  cmfb_0
timestamp 1698789667
transform 1 0 -8 0 1 -923
box 203 439 3639 2056
use integrator_new1  integrator_new1_0
timestamp 1698861456
transform 1 0 -1633 0 1 -3755
box 1247 259 5636 3705
<< end >>
