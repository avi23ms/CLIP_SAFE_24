magic
tech sky130A
magscale 1 2
timestamp 1697724144
<< nwell >>
rect -390 350 1840 1130
<< nmos >>
rect -150 -40 -120 170
rect -20 -40 10 170
rect 110 -40 140 170
rect 240 -40 270 170
rect 370 -40 400 170
rect 500 -40 530 170
rect 630 -40 660 170
rect 1010 -40 1040 170
rect 1140 -40 1170 170
rect 1270 -40 1300 170
rect 1400 -40 1430 170
rect 1530 -40 1560 170
rect 1660 -40 1690 170
<< pmos >>
rect -150 460 -120 1090
rect -20 460 10 1090
rect 110 460 140 1090
rect 240 460 270 1090
rect 370 460 400 1090
rect 500 460 530 1090
rect 630 460 660 1090
rect 1010 410 1040 1040
rect 1140 410 1170 1040
rect 1270 410 1300 1040
rect 1400 410 1430 1040
rect 1530 410 1560 1040
rect 1660 410 1690 1040
<< ndiff >>
rect -250 140 -150 170
rect -250 -10 -220 140
rect -180 -10 -150 140
rect -250 -40 -150 -10
rect -120 140 -20 170
rect -120 -10 -90 140
rect -50 -10 -20 140
rect -120 -40 -20 -10
rect 10 140 110 170
rect 10 -10 40 140
rect 80 -10 110 140
rect 10 -40 110 -10
rect 140 140 240 170
rect 140 -10 170 140
rect 210 -10 240 140
rect 140 -40 240 -10
rect 270 140 370 170
rect 270 -10 300 140
rect 340 -10 370 140
rect 270 -40 370 -10
rect 400 140 500 170
rect 400 -10 430 140
rect 470 -10 500 140
rect 400 -40 500 -10
rect 530 140 630 170
rect 530 -10 560 140
rect 600 -10 630 140
rect 530 -40 630 -10
rect 660 140 760 170
rect 660 -10 690 140
rect 730 -10 760 140
rect 660 -40 760 -10
rect 920 140 1010 170
rect 920 -10 940 140
rect 980 -10 1010 140
rect 920 -40 1010 -10
rect 1040 140 1140 170
rect 1040 -10 1070 140
rect 1110 -10 1140 140
rect 1040 -40 1140 -10
rect 1170 140 1270 170
rect 1170 -10 1200 140
rect 1240 -10 1270 140
rect 1170 -40 1270 -10
rect 1300 140 1400 170
rect 1300 -10 1330 140
rect 1370 -10 1400 140
rect 1300 -40 1400 -10
rect 1430 140 1530 170
rect 1430 -10 1460 140
rect 1500 -10 1530 140
rect 1430 -40 1530 -10
rect 1560 140 1660 170
rect 1560 -10 1590 140
rect 1630 -10 1660 140
rect 1560 -40 1660 -10
rect 1690 140 1790 170
rect 1690 -10 1720 140
rect 1760 -10 1790 140
rect 1690 -40 1790 -10
<< pdiff >>
rect -250 640 -150 1090
rect -250 490 -220 640
rect -180 490 -150 640
rect -250 460 -150 490
rect -120 1060 -20 1090
rect -120 490 -90 1060
rect -50 490 -20 1060
rect -120 460 -20 490
rect 10 1060 110 1090
rect 10 490 40 1060
rect 80 490 110 1060
rect 10 460 110 490
rect 140 1060 240 1090
rect 140 490 170 1060
rect 210 490 240 1060
rect 140 460 240 490
rect 270 1060 370 1090
rect 270 490 300 1060
rect 340 490 370 1060
rect 270 460 370 490
rect 400 1060 500 1090
rect 400 490 430 1060
rect 470 490 500 1060
rect 400 460 500 490
rect 530 1060 630 1090
rect 530 490 560 1060
rect 600 490 630 1060
rect 530 460 630 490
rect 660 1060 760 1090
rect 660 490 690 1060
rect 730 490 760 1060
rect 660 460 760 490
rect 920 1010 1010 1040
rect 920 440 940 1010
rect 980 440 1010 1010
rect 920 410 1010 440
rect 1040 1010 1140 1040
rect 1040 440 1070 1010
rect 1110 440 1140 1010
rect 1040 410 1140 440
rect 1170 1010 1270 1040
rect 1170 440 1200 1010
rect 1240 440 1270 1010
rect 1170 410 1270 440
rect 1300 1010 1400 1040
rect 1300 440 1330 1010
rect 1370 440 1400 1010
rect 1300 410 1400 440
rect 1430 1010 1530 1040
rect 1430 440 1460 1010
rect 1500 440 1530 1010
rect 1430 410 1530 440
rect 1560 1010 1660 1040
rect 1560 440 1590 1010
rect 1630 440 1660 1010
rect 1560 410 1660 440
rect 1690 1010 1790 1040
rect 1690 440 1720 1010
rect 1760 440 1790 1010
rect 1690 410 1790 440
<< ndiffc >>
rect -220 -10 -180 140
rect -90 -10 -50 140
rect 40 -10 80 140
rect 170 -10 210 140
rect 300 -10 340 140
rect 430 -10 470 140
rect 560 -10 600 140
rect 690 -10 730 140
rect 940 -10 980 140
rect 1070 -10 1110 140
rect 1200 -10 1240 140
rect 1330 -10 1370 140
rect 1460 -10 1500 140
rect 1590 -10 1630 140
rect 1720 -10 1760 140
<< pdiffc >>
rect -220 490 -180 640
rect -90 490 -50 1060
rect 40 490 80 1060
rect 170 490 210 1060
rect 300 490 340 1060
rect 430 490 470 1060
rect 560 490 600 1060
rect 690 490 730 1060
rect 940 440 980 1010
rect 1070 440 1110 1010
rect 1200 440 1240 1010
rect 1330 440 1370 1010
rect 1460 440 1500 1010
rect 1590 440 1630 1010
rect 1720 440 1760 1010
<< psubdiff >>
rect -410 140 -310 170
rect -410 -10 -380 140
rect -340 -10 -310 140
rect -410 -40 -310 -10
rect 830 140 920 170
rect 830 -10 860 140
rect 900 -10 920 140
rect 830 -40 920 -10
<< nsubdiff >>
rect -350 640 -250 1090
rect -350 490 -320 640
rect -270 490 -250 640
rect -350 460 -250 490
rect 830 1010 920 1040
rect 830 440 860 1010
rect 900 440 920 1010
rect 830 410 920 440
<< psubdiffcont >>
rect -380 -10 -340 140
rect 860 -10 900 140
<< nsubdiffcont >>
rect -320 490 -270 640
rect 860 440 900 1010
<< poly >>
rect -150 1090 -120 1120
rect -20 1110 660 1140
rect -20 1090 10 1110
rect 110 1090 140 1110
rect 240 1090 270 1110
rect 370 1090 400 1110
rect 500 1090 530 1110
rect 630 1090 660 1110
rect 1010 1040 1040 1070
rect 1140 1040 1170 1070
rect 1270 1040 1300 1070
rect 1400 1040 1430 1070
rect 1530 1040 1560 1070
rect 1660 1040 1690 1070
rect -150 170 -120 460
rect -20 440 10 460
rect 110 440 140 460
rect 240 440 270 460
rect 370 440 400 460
rect 500 440 530 460
rect 630 440 660 460
rect -20 410 660 440
rect -20 220 10 410
rect 1010 390 1040 410
rect 1140 390 1170 410
rect 1270 390 1300 410
rect 1400 390 1430 410
rect 1530 390 1560 410
rect 1660 390 1690 410
rect 1010 360 1690 390
rect 1010 340 1040 360
rect 840 320 1040 340
rect 840 270 860 320
rect 910 270 1040 320
rect 840 250 1040 270
rect 1010 220 1040 250
rect -20 190 660 220
rect -20 170 10 190
rect 110 170 140 190
rect 240 170 270 190
rect 370 170 400 190
rect 500 170 530 190
rect 630 170 660 190
rect 1010 190 1690 220
rect 1010 170 1040 190
rect 1140 170 1170 190
rect 1270 170 1300 190
rect 1400 170 1430 190
rect 1530 170 1560 190
rect 1660 170 1690 190
rect -150 -80 -120 -40
rect -20 -60 10 -40
rect 110 -60 140 -40
rect 240 -60 270 -40
rect 370 -60 400 -40
rect 500 -60 530 -40
rect 630 -60 660 -40
rect -20 -90 660 -60
rect 1010 -60 1040 -40
rect 1140 -60 1170 -40
rect 1270 -60 1300 -40
rect 1400 -60 1430 -40
rect 1530 -60 1560 -40
rect 1660 -60 1690 -40
rect 1010 -90 1690 -60
<< polycont >>
rect 860 270 910 320
<< locali >>
rect -340 1060 -160 1080
rect -340 490 -320 1060
rect -270 640 -160 1060
rect -270 490 -220 640
rect -180 490 -160 640
rect -340 470 -160 490
rect -110 1060 -30 1080
rect -110 490 -90 1060
rect -50 490 -30 1060
rect -110 470 -30 490
rect 20 1060 100 1080
rect 20 490 40 1060
rect 80 490 100 1060
rect 20 470 100 490
rect 150 1060 230 1090
rect 150 490 170 1060
rect 210 490 230 1060
rect 150 470 230 490
rect 280 1060 360 1080
rect 280 490 300 1060
rect 340 490 360 1060
rect 280 470 360 490
rect 410 1060 490 1080
rect 410 490 430 1060
rect 470 490 490 1060
rect 410 470 490 490
rect 540 1060 620 1080
rect 540 490 560 1060
rect 600 490 620 1060
rect 540 470 620 490
rect 670 1060 750 1080
rect 670 490 690 1060
rect 730 490 750 1060
rect 670 470 750 490
rect 840 1010 1000 1030
rect 840 440 860 1010
rect 900 440 940 1010
rect 980 440 1000 1010
rect 840 420 1000 440
rect 1050 1010 1130 1030
rect 1050 440 1070 1010
rect 1110 440 1130 1010
rect 1050 420 1130 440
rect 1180 1010 1260 1030
rect 1180 440 1200 1010
rect 1240 440 1260 1010
rect 1180 420 1260 440
rect 1310 1010 1390 1030
rect 1310 440 1330 1010
rect 1370 440 1390 1010
rect 1310 420 1390 440
rect 1440 1010 1520 1030
rect 1440 440 1460 1010
rect 1500 440 1520 1010
rect 1440 420 1520 440
rect 1570 1010 1650 1030
rect 1570 440 1590 1010
rect 1630 440 1650 1010
rect 1570 420 1650 440
rect 1700 1010 1780 1030
rect 1700 440 1720 1010
rect 1760 440 1780 1010
rect 1700 420 1780 440
rect 790 320 940 340
rect 790 270 860 320
rect 910 270 940 320
rect 790 250 940 270
rect -400 140 -320 160
rect -400 -10 -380 140
rect -340 -10 -320 140
rect -400 -30 -320 -10
rect -240 140 -160 160
rect -240 -10 -220 140
rect -180 -10 -160 140
rect -240 -30 -160 -10
rect -110 140 -30 160
rect -110 -10 -90 140
rect -50 -10 -30 140
rect -110 -30 -30 -10
rect 20 140 100 160
rect 20 -10 40 140
rect 80 -10 100 140
rect 20 -30 100 -10
rect 150 140 230 160
rect 150 -10 170 140
rect 210 -10 230 140
rect 150 -30 230 -10
rect 280 140 360 160
rect 280 -10 300 140
rect 340 -10 360 140
rect 280 -30 360 -10
rect 410 140 490 160
rect 410 -10 430 140
rect 470 -10 490 140
rect 410 -30 490 -10
rect 540 140 620 160
rect 540 -10 560 140
rect 600 -10 620 140
rect 540 -30 620 -10
rect 670 140 750 160
rect 670 -10 690 140
rect 730 -10 750 140
rect 670 -30 750 -10
rect 840 140 1000 160
rect 840 -10 860 140
rect 900 -10 940 140
rect 980 -10 1000 140
rect 840 -30 1000 -10
rect 1050 140 1130 160
rect 1050 -10 1070 140
rect 1110 -10 1130 140
rect 1050 -30 1130 -10
rect 1180 140 1260 160
rect 1180 -10 1200 140
rect 1240 -10 1260 140
rect 1180 -30 1260 -10
rect 1310 140 1390 160
rect 1310 -10 1330 140
rect 1370 -10 1390 140
rect 1310 -30 1390 -10
rect 1440 140 1520 160
rect 1440 -10 1460 140
rect 1500 -10 1520 140
rect 1440 -30 1520 -10
rect 1570 140 1650 160
rect 1570 -10 1590 140
rect 1630 -10 1650 140
rect 1570 -30 1650 -10
rect 1700 140 1780 160
rect 1700 -10 1720 140
rect 1760 -10 1780 140
rect 1700 -30 1780 -10
<< viali >>
rect -320 640 -270 1060
rect -320 490 -270 640
rect -90 490 -50 1060
rect 40 490 80 1060
rect 170 490 210 1060
rect 300 490 340 1060
rect 430 490 470 1060
rect 560 490 600 1060
rect 690 490 730 1060
rect 860 440 900 1010
rect 1070 440 1110 1010
rect 1200 440 1240 1010
rect 1330 440 1370 1010
rect 1460 440 1500 1010
rect 1590 440 1630 1010
rect 1720 440 1760 1010
rect 860 270 910 320
rect -380 -10 -340 140
rect -220 -10 -180 140
rect -90 -10 -50 140
rect 40 -10 80 140
rect 170 -10 210 140
rect 300 -10 340 140
rect 430 -10 470 140
rect 560 -10 600 140
rect 690 -10 730 140
rect 860 -10 900 140
rect 1070 -10 1110 140
rect 1200 -10 1240 140
rect 1330 -10 1370 140
rect 1460 -10 1500 140
rect 1590 -10 1630 140
rect 1720 -10 1760 140
<< metal1 >>
rect -340 1150 1780 1190
rect -340 1060 -260 1150
rect -340 490 -320 1060
rect -270 490 -260 1060
rect -340 470 -260 490
rect -110 1060 -30 1080
rect -110 490 -90 1060
rect -50 490 -30 1060
rect -110 340 -30 490
rect 20 1060 100 1150
rect 20 490 40 1060
rect 80 490 100 1060
rect 20 470 100 490
rect 150 1060 230 1080
rect 150 490 170 1060
rect 210 490 230 1060
rect 150 340 230 490
rect 280 1060 360 1150
rect 280 490 300 1060
rect 340 490 360 1060
rect 280 470 360 490
rect 410 1060 490 1080
rect 410 490 430 1060
rect 470 490 490 1060
rect 410 340 490 490
rect 540 1060 620 1150
rect 840 1140 1780 1150
rect 540 490 560 1060
rect 600 490 620 1060
rect 540 470 620 490
rect 670 1060 750 1080
rect 670 490 690 1060
rect 730 490 750 1060
rect 670 340 750 490
rect 840 1010 910 1140
rect 840 440 860 1010
rect 900 440 910 1010
rect 840 420 910 440
rect 1050 1010 1130 1050
rect 1050 440 1070 1010
rect 1110 440 1130 1010
rect 1050 340 1130 440
rect 1180 1010 1260 1140
rect 1180 440 1200 1010
rect 1240 440 1260 1010
rect 1180 420 1260 440
rect 1310 1010 1390 1050
rect 1310 440 1330 1010
rect 1370 440 1390 1010
rect 1310 340 1390 440
rect 1440 1010 1520 1140
rect 1440 440 1460 1010
rect 1500 440 1520 1010
rect 1440 420 1520 440
rect 1570 1010 1650 1050
rect 1570 440 1590 1010
rect 1630 440 1650 1010
rect 1570 340 1650 440
rect 1700 1010 1780 1140
rect 1700 440 1720 1010
rect 1760 440 1780 1010
rect 1700 420 1780 440
rect -240 320 980 340
rect -240 310 860 320
rect -400 140 -320 160
rect -400 -10 -380 140
rect -340 -10 -320 140
rect -400 -100 -320 -10
rect -240 140 -160 310
rect 790 270 860 310
rect 910 270 980 320
rect -240 -10 -220 140
rect -180 -10 -160 140
rect -240 -30 -160 -10
rect -110 230 750 260
rect 790 250 980 270
rect 1050 300 1650 340
rect -110 140 -30 230
rect 150 200 230 230
rect -110 -10 -90 140
rect -50 -10 -30 140
rect 0 140 230 200
rect 0 0 40 140
rect -110 -30 -30 -10
rect 20 -10 40 0
rect 80 0 170 140
rect 80 -10 100 0
rect 20 -100 100 -10
rect 150 -10 170 0
rect 210 -10 230 140
rect 150 -30 230 -10
rect 280 140 360 160
rect 280 -10 300 140
rect 340 -10 360 140
rect 280 -100 360 -10
rect 410 140 490 230
rect 410 -10 430 140
rect 470 -10 490 140
rect 410 -30 490 -10
rect 540 140 620 160
rect 540 -10 560 140
rect 600 -10 620 140
rect 540 -100 620 -10
rect 670 140 750 230
rect 670 -10 690 140
rect 730 -10 750 140
rect 670 -20 750 -10
rect 840 140 910 160
rect 840 -10 860 140
rect 900 -10 910 140
rect 840 -100 910 -10
rect 1050 140 1130 300
rect 1050 -10 1070 140
rect 1110 -10 1130 140
rect 1050 -30 1130 -10
rect 1180 140 1260 160
rect 1180 -10 1200 140
rect 1240 -10 1260 140
rect 1180 -100 1260 -10
rect 1310 140 1390 300
rect 1310 -10 1330 140
rect 1370 -10 1390 140
rect 1310 -30 1390 -10
rect 1440 140 1520 160
rect 1440 -10 1460 140
rect 1500 -10 1520 140
rect 1440 -100 1520 -10
rect 1570 140 1650 300
rect 1570 -10 1590 140
rect 1630 -10 1650 140
rect 1570 -30 1650 -10
rect 1700 140 1780 160
rect 1700 -10 1720 140
rect 1760 -10 1780 140
rect 1700 -100 1780 -10
rect -400 -130 1780 -100
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__pfet_01v8_XGSNAL  XM1
timestamp 0
transform 1 0 527 0 1 1013
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_XGSNAL  XM2
timestamp 0
transform 1 0 158 0 1 1066
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_ATLS57  XM4
timestamp 0
transform 1 0 896 0 1 851
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_ATLS57  XM5
timestamp 0
transform 1 0 1265 0 1 798
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 GND
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 B
port 4 nsew
<< end >>
