magic
tech sky130A
timestamp 1698622134
<< error_p >>
rect -277 57 -248 60
rect -67 57 -38 60
rect 143 57 172 60
rect 353 57 382 60
rect -277 40 -271 57
rect -67 40 -61 57
rect 143 40 149 57
rect 353 40 359 57
rect -277 37 -248 40
rect -67 37 -38 40
rect 143 37 172 40
rect 353 37 382 40
rect -382 -40 -353 -37
rect -172 -40 -143 -37
rect 38 -40 67 -37
rect 248 -40 277 -37
rect -382 -57 -376 -40
rect -172 -57 -166 -40
rect 38 -57 44 -40
rect 248 -57 254 -40
rect -382 -60 -353 -57
rect -172 -60 -143 -57
rect 38 -60 67 -57
rect 248 -60 277 -57
<< nmos >>
rect -375 -21 -360 21
rect -270 -21 -255 21
rect -165 -21 -150 21
rect -60 -21 -45 21
rect 45 -21 60 21
rect 150 -21 165 21
rect 255 -21 270 21
rect 360 -21 375 21
<< ndiff >>
rect -406 15 -375 21
rect -406 -15 -400 15
rect -383 -15 -375 15
rect -406 -21 -375 -15
rect -360 15 -329 21
rect -360 -15 -352 15
rect -335 -15 -329 15
rect -360 -21 -329 -15
rect -301 15 -270 21
rect -301 -15 -295 15
rect -278 -15 -270 15
rect -301 -21 -270 -15
rect -255 15 -224 21
rect -255 -15 -247 15
rect -230 -15 -224 15
rect -255 -21 -224 -15
rect -196 15 -165 21
rect -196 -15 -190 15
rect -173 -15 -165 15
rect -196 -21 -165 -15
rect -150 15 -119 21
rect -150 -15 -142 15
rect -125 -15 -119 15
rect -150 -21 -119 -15
rect -91 15 -60 21
rect -91 -15 -85 15
rect -68 -15 -60 15
rect -91 -21 -60 -15
rect -45 15 -14 21
rect -45 -15 -37 15
rect -20 -15 -14 15
rect -45 -21 -14 -15
rect 14 15 45 21
rect 14 -15 20 15
rect 37 -15 45 15
rect 14 -21 45 -15
rect 60 15 91 21
rect 60 -15 68 15
rect 85 -15 91 15
rect 60 -21 91 -15
rect 119 15 150 21
rect 119 -15 125 15
rect 142 -15 150 15
rect 119 -21 150 -15
rect 165 15 196 21
rect 165 -15 173 15
rect 190 -15 196 15
rect 165 -21 196 -15
rect 224 15 255 21
rect 224 -15 230 15
rect 247 -15 255 15
rect 224 -21 255 -15
rect 270 15 301 21
rect 270 -15 278 15
rect 295 -15 301 15
rect 270 -21 301 -15
rect 329 15 360 21
rect 329 -15 335 15
rect 352 -15 360 15
rect 329 -21 360 -15
rect 375 15 406 21
rect 375 -15 383 15
rect 400 -15 406 15
rect 375 -21 406 -15
<< ndiffc >>
rect -400 -15 -383 15
rect -352 -15 -335 15
rect -295 -15 -278 15
rect -247 -15 -230 15
rect -190 -15 -173 15
rect -142 -15 -125 15
rect -85 -15 -68 15
rect -37 -15 -20 15
rect 20 -15 37 15
rect 68 -15 85 15
rect 125 -15 142 15
rect 173 -15 190 15
rect 230 -15 247 15
rect 278 -15 295 15
rect 335 -15 352 15
rect 383 -15 400 15
<< poly >>
rect -279 57 -246 65
rect -279 40 -271 57
rect -254 40 -246 57
rect -375 21 -360 34
rect -279 32 -246 40
rect -69 57 -36 65
rect -69 40 -61 57
rect -44 40 -36 57
rect -270 21 -255 32
rect -165 21 -150 34
rect -69 32 -36 40
rect 141 57 174 65
rect 141 40 149 57
rect 166 40 174 57
rect -60 21 -45 32
rect 45 21 60 34
rect 141 32 174 40
rect 351 57 384 65
rect 351 40 359 57
rect 376 40 384 57
rect 150 21 165 32
rect 255 21 270 34
rect 351 32 384 40
rect 360 21 375 32
rect -375 -32 -360 -21
rect -384 -40 -351 -32
rect -270 -34 -255 -21
rect -165 -32 -150 -21
rect -384 -57 -376 -40
rect -359 -57 -351 -40
rect -384 -65 -351 -57
rect -174 -40 -141 -32
rect -60 -34 -45 -21
rect 45 -32 60 -21
rect -174 -57 -166 -40
rect -149 -57 -141 -40
rect -174 -65 -141 -57
rect 36 -40 69 -32
rect 150 -34 165 -21
rect 255 -32 270 -21
rect 36 -57 44 -40
rect 61 -57 69 -40
rect 36 -65 69 -57
rect 246 -40 279 -32
rect 360 -34 375 -21
rect 246 -57 254 -40
rect 271 -57 279 -40
rect 246 -65 279 -57
<< polycont >>
rect -271 40 -254 57
rect -61 40 -44 57
rect 149 40 166 57
rect 359 40 376 57
rect -376 -57 -359 -40
rect -166 -57 -149 -40
rect 44 -57 61 -40
rect 254 -57 271 -40
<< locali >>
rect -279 40 -271 57
rect -254 40 -246 57
rect -69 40 -61 57
rect -44 40 -36 57
rect 141 40 149 57
rect 166 40 174 57
rect 351 40 359 57
rect 376 40 384 57
rect -400 15 -383 23
rect -400 -23 -383 -15
rect -352 15 -335 23
rect -352 -23 -335 -15
rect -295 15 -278 23
rect -295 -23 -278 -15
rect -247 15 -230 23
rect -247 -23 -230 -15
rect -190 15 -173 23
rect -190 -23 -173 -15
rect -142 15 -125 23
rect -142 -23 -125 -15
rect -85 15 -68 23
rect -85 -23 -68 -15
rect -37 15 -20 23
rect -37 -23 -20 -15
rect 20 15 37 23
rect 20 -23 37 -15
rect 68 15 85 23
rect 68 -23 85 -15
rect 125 15 142 23
rect 125 -23 142 -15
rect 173 15 190 23
rect 173 -23 190 -15
rect 230 15 247 23
rect 230 -23 247 -15
rect 278 15 295 23
rect 278 -23 295 -15
rect 335 15 352 23
rect 335 -23 352 -15
rect 383 15 400 23
rect 383 -23 400 -15
rect -384 -57 -376 -40
rect -359 -57 -351 -40
rect -174 -57 -166 -40
rect -149 -57 -141 -40
rect 36 -57 44 -40
rect 61 -57 69 -40
rect 246 -57 254 -40
rect 271 -57 279 -40
<< viali >>
rect -271 40 -254 57
rect -61 40 -44 57
rect 149 40 166 57
rect 359 40 376 57
rect -400 -15 -383 15
rect -352 -15 -335 15
rect -295 -15 -278 15
rect -247 -15 -230 15
rect -190 -15 -173 15
rect -142 -15 -125 15
rect -85 -15 -68 15
rect -37 -15 -20 15
rect 20 -15 37 15
rect 68 -15 85 15
rect 125 -15 142 15
rect 173 -15 190 15
rect 230 -15 247 15
rect 278 -15 295 15
rect 335 -15 352 15
rect 383 -15 400 15
rect -376 -57 -359 -40
rect -166 -57 -149 -40
rect 44 -57 61 -40
rect 254 -57 271 -40
<< metal1 >>
rect -277 57 -248 60
rect -277 40 -271 57
rect -254 40 -248 57
rect -277 37 -248 40
rect -67 57 -38 60
rect -67 40 -61 57
rect -44 40 -38 57
rect -67 37 -38 40
rect 143 57 172 60
rect 143 40 149 57
rect 166 40 172 57
rect 143 37 172 40
rect 353 57 382 60
rect 353 40 359 57
rect 376 40 382 57
rect 353 37 382 40
rect -403 15 -380 21
rect -403 -15 -400 15
rect -383 -15 -380 15
rect -403 -21 -380 -15
rect -355 15 -332 21
rect -355 -15 -352 15
rect -335 -15 -332 15
rect -355 -21 -332 -15
rect -298 15 -275 21
rect -298 -15 -295 15
rect -278 -15 -275 15
rect -298 -21 -275 -15
rect -250 15 -227 21
rect -250 -15 -247 15
rect -230 -15 -227 15
rect -250 -21 -227 -15
rect -193 15 -170 21
rect -193 -15 -190 15
rect -173 -15 -170 15
rect -193 -21 -170 -15
rect -145 15 -122 21
rect -145 -15 -142 15
rect -125 -15 -122 15
rect -145 -21 -122 -15
rect -88 15 -65 21
rect -88 -15 -85 15
rect -68 -15 -65 15
rect -88 -21 -65 -15
rect -40 15 -17 21
rect -40 -15 -37 15
rect -20 -15 -17 15
rect -40 -21 -17 -15
rect 17 15 40 21
rect 17 -15 20 15
rect 37 -15 40 15
rect 17 -21 40 -15
rect 65 15 88 21
rect 65 -15 68 15
rect 85 -15 88 15
rect 65 -21 88 -15
rect 122 15 145 21
rect 122 -15 125 15
rect 142 -15 145 15
rect 122 -21 145 -15
rect 170 15 193 21
rect 170 -15 173 15
rect 190 -15 193 15
rect 170 -21 193 -15
rect 227 15 250 21
rect 227 -15 230 15
rect 247 -15 250 15
rect 227 -21 250 -15
rect 275 15 298 21
rect 275 -15 278 15
rect 295 -15 298 15
rect 275 -21 298 -15
rect 332 15 355 21
rect 332 -15 335 15
rect 352 -15 355 15
rect 332 -21 355 -15
rect 380 15 403 21
rect 380 -15 383 15
rect 400 -15 403 15
rect 380 -21 403 -15
rect -382 -40 -353 -37
rect -382 -57 -376 -40
rect -359 -57 -353 -40
rect -382 -60 -353 -57
rect -172 -40 -143 -37
rect -172 -57 -166 -40
rect -149 -57 -143 -40
rect -172 -60 -143 -57
rect 38 -40 67 -37
rect 38 -57 44 -40
rect 61 -57 67 -40
rect 38 -60 67 -57
rect 248 -40 277 -37
rect 248 -57 254 -40
rect 271 -57 277 -40
rect 248 -60 277 -57
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
