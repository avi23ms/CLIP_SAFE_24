magic
tech sky130A
magscale 1 2
timestamp 1698771642
<< locali >>
rect 30 2142 2584 2181
rect 30 2103 89 2142
rect 30 2070 2584 2103
rect 169 1755 316 1838
rect 554 1748 700 1814
rect 1980 1736 2134 1834
rect 2367 1752 2521 1830
rect 179 1135 319 1212
rect 554 1135 702 1210
rect 1984 1128 2138 1206
rect 2369 1137 2523 1215
rect 238 913 2674 951
rect 238 874 260 913
rect 2656 874 2674 913
rect 238 840 2674 874
<< viali >>
rect 89 2103 2584 2142
rect 260 874 2656 913
<< metal1 >>
rect 30 2148 2584 2181
rect 30 2142 2596 2148
rect 30 2103 89 2142
rect 2584 2103 2596 2142
rect 30 2097 2596 2103
rect 30 2070 2584 2097
rect 330 1963 340 2020
rect 409 1963 419 2020
rect 724 1961 734 2018
rect 803 1961 813 2018
rect 334 1315 344 1372
rect 413 1315 423 1372
rect 454 1219 491 1918
rect 822 1732 1090 1908
rect 1128 1687 1163 2004
rect 722 1630 732 1687
rect 801 1630 811 1687
rect 1100 1630 1110 1687
rect 1189 1630 1199 1687
rect 1128 1379 1163 1630
rect 1097 1325 1107 1379
rect 1182 1325 1192 1379
rect 432 1167 442 1219
rect 430 1104 440 1167
rect 496 1156 506 1219
rect 494 1104 504 1156
rect 454 1098 491 1104
rect 827 1096 1095 1272
rect 716 998 726 1055
rect 795 998 805 1055
rect 1128 1051 1163 1325
rect 1228 1255 1261 1910
rect 1212 1200 1222 1255
rect 1279 1200 1289 1255
rect 1427 1201 1460 1916
rect 1515 1380 1550 2004
rect 1878 1968 1975 2022
rect 2260 1962 2270 2018
rect 2374 1962 2384 2018
rect 1601 1730 1869 1906
rect 2195 1874 2232 1916
rect 2186 1817 2196 1874
rect 2182 1750 2192 1817
rect 2255 1807 2265 1874
rect 2251 1750 2261 1807
rect 1858 1624 1868 1680
rect 1972 1624 1982 1680
rect 1501 1323 1511 1380
rect 1589 1323 1599 1380
rect 1228 1161 1261 1200
rect 1208 1106 1218 1161
rect 1275 1106 1285 1161
rect 1388 1147 1398 1201
rect 1473 1150 1483 1201
rect 1228 1090 1261 1106
rect 1390 1096 1400 1147
rect 1475 1096 1485 1150
rect 1515 1052 1550 1323
rect 1884 1315 1981 1369
rect 1595 1096 1863 1272
rect 2195 1096 2232 1750
rect 2266 1626 2363 1680
rect 2272 1369 2282 1376
rect 2268 1320 2282 1369
rect 2386 1320 2396 1376
rect 2268 1315 2365 1320
rect 1108 997 1118 1051
rect 1193 997 1203 1051
rect 1505 995 1515 1052
rect 1593 995 1603 1052
rect 1878 998 1888 1054
rect 1992 998 2002 1054
rect 238 913 2674 951
rect 238 874 260 913
rect 2656 874 2674 913
rect 238 840 2674 874
<< via1 >>
rect 340 1963 409 2020
rect 734 1961 803 2018
rect 344 1315 413 1372
rect 732 1630 801 1687
rect 1110 1630 1189 1687
rect 1107 1325 1182 1379
rect 442 1167 496 1219
rect 440 1156 496 1167
rect 440 1104 494 1156
rect 726 998 795 1055
rect 1222 1200 1279 1255
rect 2270 1962 2374 2018
rect 2196 1817 2255 1874
rect 2192 1807 2255 1817
rect 2192 1750 2251 1807
rect 1868 1624 1972 1680
rect 1511 1323 1589 1380
rect 1218 1106 1275 1161
rect 1398 1150 1473 1201
rect 1398 1147 1475 1150
rect 1400 1096 1475 1147
rect 2282 1320 2386 1376
rect 1118 997 1193 1051
rect 1515 995 1593 1052
rect 1888 998 1992 1054
<< metal2 >>
rect 2284 2078 2512 2110
rect 340 2020 409 2030
rect 2284 2028 2316 2078
rect 171 1967 340 2006
rect 171 917 210 1967
rect 340 1953 409 1963
rect 734 2018 803 2028
rect 734 1951 803 1961
rect 2270 2018 2374 2028
rect 2270 1952 2374 1962
rect 2196 1874 2255 1884
rect 1133 1817 2196 1827
rect 1133 1771 2192 1817
rect 1133 1697 1189 1771
rect 2251 1797 2255 1807
rect 2192 1740 2251 1750
rect 732 1687 801 1697
rect 732 1620 801 1630
rect 1110 1687 1189 1697
rect 1110 1620 1189 1630
rect 1868 1680 1972 1690
rect 742 1592 781 1620
rect 1868 1614 1972 1624
rect 742 1572 780 1592
rect 341 1534 780 1572
rect 1898 1581 1932 1614
rect 1898 1547 2319 1581
rect 341 1382 379 1534
rect 1898 1532 1932 1547
rect 455 1467 1557 1498
rect 455 1411 486 1467
rect 1229 1411 1260 1467
rect 1526 1411 1557 1467
rect 341 1372 413 1382
rect 341 1315 344 1372
rect 341 1305 413 1315
rect 450 1378 486 1411
rect 1107 1379 1182 1411
rect 341 1302 379 1305
rect 450 1229 485 1378
rect 1107 1315 1182 1325
rect 442 1219 496 1229
rect 440 1167 442 1177
rect 494 1146 496 1156
rect 440 1094 494 1104
rect 726 1055 795 1065
rect 1139 1061 1173 1315
rect 1224 1265 1260 1411
rect 1511 1390 1557 1411
rect 1511 1380 1589 1390
rect 2285 1386 2319 1547
rect 1511 1313 1589 1323
rect 2282 1376 2386 1386
rect 1222 1255 1279 1265
rect 1216 1200 1222 1212
rect 1279 1200 1281 1212
rect 1216 1161 1281 1200
rect 1216 1137 1218 1161
rect 1275 1137 1281 1161
rect 1398 1201 1473 1211
rect 1473 1150 1475 1160
rect 1398 1137 1400 1147
rect 1218 1096 1275 1106
rect 1400 1086 1475 1096
rect 726 988 795 998
rect 1118 1053 1193 1061
rect 1433 1053 1467 1086
rect 1526 1062 1557 1313
rect 2282 1310 2386 1320
rect 1118 1051 1467 1053
rect 1193 1019 1467 1051
rect 1433 1018 1467 1019
rect 1515 1052 1593 1062
rect 747 917 786 988
rect 1118 987 1193 997
rect 1515 985 1593 995
rect 1888 1054 1992 1064
rect 1888 988 1992 998
rect 171 878 786 917
rect 1936 918 1968 988
rect 2480 918 2512 2078
rect 1936 886 2512 918
use sky130_fd_pr__pfet_01v8_X3YSY6  sky130_fd_pr__pfet_01v8_X3YSY6_0
timestamp 1698771642
transform 1 0 2308 0 1 1821
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_X3YSY6  XM13
timestamp 1698771642
transform 1 0 378 0 1 1821
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_X3YSY6  XM14
timestamp 1698771642
transform 1 0 764 0 1 1821
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_X3YSY6  XM15
timestamp 1698771642
transform 1 0 1150 0 1 1821
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_X3YSY6  XM16
timestamp 1698771642
transform 1 0 1536 0 1 1821
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_X3YSY6  XM17
timestamp 1698771642
transform 1 0 1922 0 1 1821
box -246 -319 246 319
use sky130_fd_pr__nfet_01v8_PVEW3M  XM19
timestamp 1698771642
transform 1 0 1924 0 1 1185
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM20
timestamp 1698771642
transform 1 0 2310 0 1 1185
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM21
timestamp 1698771642
transform 1 0 380 0 1 1185
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM22
timestamp 1698771642
transform 1 0 766 0 1 1185
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM23
timestamp 1698771642
transform 1 0 1152 0 1 1185
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_PVEW3M  XM24
timestamp 1698771642
transform 1 0 1538 0 1 1185
box -246 -310 246 310
<< end >>
