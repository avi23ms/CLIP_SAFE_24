magic
tech sky130A
magscale 1 2
timestamp 1698657458
<< nwell >>
rect -1649 104 1649 142
rect -1745 -142 1745 104
<< pmos >>
rect -1647 -42 -1617 42
rect -1551 -42 -1521 42
rect -1455 -42 -1425 42
rect -1359 -42 -1329 42
rect -1263 -42 -1233 42
rect -1167 -42 -1137 42
rect -1071 -42 -1041 42
rect -975 -42 -945 42
rect -879 -42 -849 42
rect -783 -42 -753 42
rect -687 -42 -657 42
rect -591 -42 -561 42
rect -495 -42 -465 42
rect -399 -42 -369 42
rect -303 -42 -273 42
rect -207 -42 -177 42
rect -111 -42 -81 42
rect -15 -42 15 42
rect 81 -42 111 42
rect 177 -42 207 42
rect 273 -42 303 42
rect 369 -42 399 42
rect 465 -42 495 42
rect 561 -42 591 42
rect 657 -42 687 42
rect 753 -42 783 42
rect 849 -42 879 42
rect 945 -42 975 42
rect 1041 -42 1071 42
rect 1137 -42 1167 42
rect 1233 -42 1263 42
rect 1329 -42 1359 42
rect 1425 -42 1455 42
rect 1521 -42 1551 42
rect 1617 -42 1647 42
<< pdiff >>
rect -1709 30 -1647 42
rect -1709 -30 -1697 30
rect -1663 -30 -1647 30
rect -1709 -42 -1647 -30
rect -1617 30 -1551 42
rect -1617 -30 -1601 30
rect -1567 -30 -1551 30
rect -1617 -42 -1551 -30
rect -1521 30 -1455 42
rect -1521 -30 -1505 30
rect -1471 -30 -1455 30
rect -1521 -42 -1455 -30
rect -1425 30 -1359 42
rect -1425 -30 -1409 30
rect -1375 -30 -1359 30
rect -1425 -42 -1359 -30
rect -1329 30 -1263 42
rect -1329 -30 -1313 30
rect -1279 -30 -1263 30
rect -1329 -42 -1263 -30
rect -1233 30 -1167 42
rect -1233 -30 -1217 30
rect -1183 -30 -1167 30
rect -1233 -42 -1167 -30
rect -1137 30 -1071 42
rect -1137 -30 -1121 30
rect -1087 -30 -1071 30
rect -1137 -42 -1071 -30
rect -1041 30 -975 42
rect -1041 -30 -1025 30
rect -991 -30 -975 30
rect -1041 -42 -975 -30
rect -945 30 -879 42
rect -945 -30 -929 30
rect -895 -30 -879 30
rect -945 -42 -879 -30
rect -849 30 -783 42
rect -849 -30 -833 30
rect -799 -30 -783 30
rect -849 -42 -783 -30
rect -753 30 -687 42
rect -753 -30 -737 30
rect -703 -30 -687 30
rect -753 -42 -687 -30
rect -657 30 -591 42
rect -657 -30 -641 30
rect -607 -30 -591 30
rect -657 -42 -591 -30
rect -561 30 -495 42
rect -561 -30 -545 30
rect -511 -30 -495 30
rect -561 -42 -495 -30
rect -465 30 -399 42
rect -465 -30 -449 30
rect -415 -30 -399 30
rect -465 -42 -399 -30
rect -369 30 -303 42
rect -369 -30 -353 30
rect -319 -30 -303 30
rect -369 -42 -303 -30
rect -273 30 -207 42
rect -273 -30 -257 30
rect -223 -30 -207 30
rect -273 -42 -207 -30
rect -177 30 -111 42
rect -177 -30 -161 30
rect -127 -30 -111 30
rect -177 -42 -111 -30
rect -81 30 -15 42
rect -81 -30 -65 30
rect -31 -30 -15 30
rect -81 -42 -15 -30
rect 15 30 81 42
rect 15 -30 31 30
rect 65 -30 81 30
rect 15 -42 81 -30
rect 111 30 177 42
rect 111 -30 127 30
rect 161 -30 177 30
rect 111 -42 177 -30
rect 207 30 273 42
rect 207 -30 223 30
rect 257 -30 273 30
rect 207 -42 273 -30
rect 303 30 369 42
rect 303 -30 319 30
rect 353 -30 369 30
rect 303 -42 369 -30
rect 399 30 465 42
rect 399 -30 415 30
rect 449 -30 465 30
rect 399 -42 465 -30
rect 495 30 561 42
rect 495 -30 511 30
rect 545 -30 561 30
rect 495 -42 561 -30
rect 591 30 657 42
rect 591 -30 607 30
rect 641 -30 657 30
rect 591 -42 657 -30
rect 687 30 753 42
rect 687 -30 703 30
rect 737 -30 753 30
rect 687 -42 753 -30
rect 783 30 849 42
rect 783 -30 799 30
rect 833 -30 849 30
rect 783 -42 849 -30
rect 879 30 945 42
rect 879 -30 895 30
rect 929 -30 945 30
rect 879 -42 945 -30
rect 975 30 1041 42
rect 975 -30 991 30
rect 1025 -30 1041 30
rect 975 -42 1041 -30
rect 1071 30 1137 42
rect 1071 -30 1087 30
rect 1121 -30 1137 30
rect 1071 -42 1137 -30
rect 1167 30 1233 42
rect 1167 -30 1183 30
rect 1217 -30 1233 30
rect 1167 -42 1233 -30
rect 1263 30 1329 42
rect 1263 -30 1279 30
rect 1313 -30 1329 30
rect 1263 -42 1329 -30
rect 1359 30 1425 42
rect 1359 -30 1375 30
rect 1409 -30 1425 30
rect 1359 -42 1425 -30
rect 1455 30 1521 42
rect 1455 -30 1471 30
rect 1505 -30 1521 30
rect 1455 -42 1521 -30
rect 1551 30 1617 42
rect 1551 -30 1567 30
rect 1601 -30 1617 30
rect 1551 -42 1617 -30
rect 1647 30 1709 42
rect 1647 -30 1663 30
rect 1697 -30 1709 30
rect 1647 -42 1709 -30
<< pdiffc >>
rect -1697 -30 -1663 30
rect -1601 -30 -1567 30
rect -1505 -30 -1471 30
rect -1409 -30 -1375 30
rect -1313 -30 -1279 30
rect -1217 -30 -1183 30
rect -1121 -30 -1087 30
rect -1025 -30 -991 30
rect -929 -30 -895 30
rect -833 -30 -799 30
rect -737 -30 -703 30
rect -641 -30 -607 30
rect -545 -30 -511 30
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
rect 511 -30 545 30
rect 607 -30 641 30
rect 703 -30 737 30
rect 799 -30 833 30
rect 895 -30 929 30
rect 991 -30 1025 30
rect 1087 -30 1121 30
rect 1183 -30 1217 30
rect 1279 -30 1313 30
rect 1375 -30 1409 30
rect 1471 -30 1505 30
rect 1567 -30 1601 30
rect 1663 -30 1697 30
<< poly >>
rect -1569 123 -1503 139
rect -1569 89 -1553 123
rect -1519 89 -1503 123
rect -1569 73 -1503 89
rect -1377 123 -1311 139
rect -1377 89 -1361 123
rect -1327 89 -1311 123
rect -1377 73 -1311 89
rect -1185 123 -1119 139
rect -1185 89 -1169 123
rect -1135 89 -1119 123
rect -1185 73 -1119 89
rect -993 123 -927 139
rect -993 89 -977 123
rect -943 89 -927 123
rect -993 73 -927 89
rect -801 123 -735 139
rect -801 89 -785 123
rect -751 89 -735 123
rect -801 73 -735 89
rect -609 123 -543 139
rect -609 89 -593 123
rect -559 89 -543 123
rect -609 73 -543 89
rect -417 123 -351 139
rect -417 89 -401 123
rect -367 89 -351 123
rect -417 73 -351 89
rect -225 123 -159 139
rect -225 89 -209 123
rect -175 89 -159 123
rect -225 73 -159 89
rect -33 123 33 139
rect -33 89 -17 123
rect 17 89 33 123
rect -33 73 33 89
rect 159 123 225 139
rect 159 89 175 123
rect 209 89 225 123
rect 159 73 225 89
rect 351 123 417 139
rect 351 89 367 123
rect 401 89 417 123
rect 351 73 417 89
rect 543 123 609 139
rect 543 89 559 123
rect 593 89 609 123
rect 543 73 609 89
rect 735 123 801 139
rect 735 89 751 123
rect 785 89 801 123
rect 735 73 801 89
rect 927 123 993 139
rect 927 89 943 123
rect 977 89 993 123
rect 927 73 993 89
rect 1119 123 1185 139
rect 1119 89 1135 123
rect 1169 89 1185 123
rect 1119 73 1185 89
rect 1311 123 1377 139
rect 1311 89 1327 123
rect 1361 89 1377 123
rect 1311 73 1377 89
rect 1503 123 1569 139
rect 1503 89 1519 123
rect 1553 89 1569 123
rect 1503 73 1569 89
rect -1647 42 -1617 68
rect -1551 42 -1521 73
rect -1455 42 -1425 68
rect -1359 42 -1329 73
rect -1263 42 -1233 68
rect -1167 42 -1137 73
rect -1071 42 -1041 68
rect -975 42 -945 73
rect -879 42 -849 68
rect -783 42 -753 73
rect -687 42 -657 68
rect -591 42 -561 73
rect -495 42 -465 68
rect -399 42 -369 73
rect -303 42 -273 68
rect -207 42 -177 73
rect -111 42 -81 68
rect -15 42 15 73
rect 81 42 111 68
rect 177 42 207 73
rect 273 42 303 68
rect 369 42 399 73
rect 465 42 495 68
rect 561 42 591 73
rect 657 42 687 68
rect 753 42 783 73
rect 849 42 879 68
rect 945 42 975 73
rect 1041 42 1071 68
rect 1137 42 1167 73
rect 1233 42 1263 68
rect 1329 42 1359 73
rect 1425 42 1455 68
rect 1521 42 1551 73
rect 1617 42 1647 68
rect -1647 -73 -1617 -42
rect -1551 -68 -1521 -42
rect -1455 -73 -1425 -42
rect -1359 -68 -1329 -42
rect -1263 -73 -1233 -42
rect -1167 -68 -1137 -42
rect -1071 -73 -1041 -42
rect -975 -68 -945 -42
rect -879 -73 -849 -42
rect -783 -68 -753 -42
rect -687 -73 -657 -42
rect -591 -68 -561 -42
rect -495 -73 -465 -42
rect -399 -68 -369 -42
rect -303 -73 -273 -42
rect -207 -68 -177 -42
rect -111 -73 -81 -42
rect -15 -68 15 -42
rect 81 -73 111 -42
rect 177 -68 207 -42
rect 273 -73 303 -42
rect 369 -68 399 -42
rect 465 -73 495 -42
rect 561 -68 591 -42
rect 657 -73 687 -42
rect 753 -68 783 -42
rect 849 -73 879 -42
rect 945 -68 975 -42
rect 1041 -73 1071 -42
rect 1137 -68 1167 -42
rect 1233 -73 1263 -42
rect 1329 -68 1359 -42
rect 1425 -73 1455 -42
rect 1521 -68 1551 -42
rect 1617 -73 1647 -42
rect -1665 -89 -1599 -73
rect -1665 -123 -1649 -89
rect -1615 -123 -1599 -89
rect -1665 -139 -1599 -123
rect -1473 -89 -1407 -73
rect -1473 -123 -1457 -89
rect -1423 -123 -1407 -89
rect -1473 -139 -1407 -123
rect -1281 -89 -1215 -73
rect -1281 -123 -1265 -89
rect -1231 -123 -1215 -89
rect -1281 -139 -1215 -123
rect -1089 -89 -1023 -73
rect -1089 -123 -1073 -89
rect -1039 -123 -1023 -89
rect -1089 -139 -1023 -123
rect -897 -89 -831 -73
rect -897 -123 -881 -89
rect -847 -123 -831 -89
rect -897 -139 -831 -123
rect -705 -89 -639 -73
rect -705 -123 -689 -89
rect -655 -123 -639 -89
rect -705 -139 -639 -123
rect -513 -89 -447 -73
rect -513 -123 -497 -89
rect -463 -123 -447 -89
rect -513 -139 -447 -123
rect -321 -89 -255 -73
rect -321 -123 -305 -89
rect -271 -123 -255 -89
rect -321 -139 -255 -123
rect -129 -89 -63 -73
rect -129 -123 -113 -89
rect -79 -123 -63 -89
rect -129 -139 -63 -123
rect 63 -89 129 -73
rect 63 -123 79 -89
rect 113 -123 129 -89
rect 63 -139 129 -123
rect 255 -89 321 -73
rect 255 -123 271 -89
rect 305 -123 321 -89
rect 255 -139 321 -123
rect 447 -89 513 -73
rect 447 -123 463 -89
rect 497 -123 513 -89
rect 447 -139 513 -123
rect 639 -89 705 -73
rect 639 -123 655 -89
rect 689 -123 705 -89
rect 639 -139 705 -123
rect 831 -89 897 -73
rect 831 -123 847 -89
rect 881 -123 897 -89
rect 831 -139 897 -123
rect 1023 -89 1089 -73
rect 1023 -123 1039 -89
rect 1073 -123 1089 -89
rect 1023 -139 1089 -123
rect 1215 -89 1281 -73
rect 1215 -123 1231 -89
rect 1265 -123 1281 -89
rect 1215 -139 1281 -123
rect 1407 -89 1473 -73
rect 1407 -123 1423 -89
rect 1457 -123 1473 -89
rect 1407 -139 1473 -123
rect 1599 -89 1665 -73
rect 1599 -123 1615 -89
rect 1649 -123 1665 -89
rect 1599 -139 1665 -123
<< polycont >>
rect -1553 89 -1519 123
rect -1361 89 -1327 123
rect -1169 89 -1135 123
rect -977 89 -943 123
rect -785 89 -751 123
rect -593 89 -559 123
rect -401 89 -367 123
rect -209 89 -175 123
rect -17 89 17 123
rect 175 89 209 123
rect 367 89 401 123
rect 559 89 593 123
rect 751 89 785 123
rect 943 89 977 123
rect 1135 89 1169 123
rect 1327 89 1361 123
rect 1519 89 1553 123
rect -1649 -123 -1615 -89
rect -1457 -123 -1423 -89
rect -1265 -123 -1231 -89
rect -1073 -123 -1039 -89
rect -881 -123 -847 -89
rect -689 -123 -655 -89
rect -497 -123 -463 -89
rect -305 -123 -271 -89
rect -113 -123 -79 -89
rect 79 -123 113 -89
rect 271 -123 305 -89
rect 463 -123 497 -89
rect 655 -123 689 -89
rect 847 -123 881 -89
rect 1039 -123 1073 -89
rect 1231 -123 1265 -89
rect 1423 -123 1457 -89
rect 1615 -123 1649 -89
<< locali >>
rect -1569 89 -1553 123
rect -1519 89 -1503 123
rect -1377 89 -1361 123
rect -1327 89 -1311 123
rect -1185 89 -1169 123
rect -1135 89 -1119 123
rect -993 89 -977 123
rect -943 89 -927 123
rect -801 89 -785 123
rect -751 89 -735 123
rect -609 89 -593 123
rect -559 89 -543 123
rect -417 89 -401 123
rect -367 89 -351 123
rect -225 89 -209 123
rect -175 89 -159 123
rect -33 89 -17 123
rect 17 89 33 123
rect 159 89 175 123
rect 209 89 225 123
rect 351 89 367 123
rect 401 89 417 123
rect 543 89 559 123
rect 593 89 609 123
rect 735 89 751 123
rect 785 89 801 123
rect 927 89 943 123
rect 977 89 993 123
rect 1119 89 1135 123
rect 1169 89 1185 123
rect 1311 89 1327 123
rect 1361 89 1377 123
rect 1503 89 1519 123
rect 1553 89 1569 123
rect -1697 30 -1663 46
rect -1697 -46 -1663 -30
rect -1601 30 -1567 46
rect -1601 -46 -1567 -30
rect -1505 30 -1471 46
rect -1505 -46 -1471 -30
rect -1409 30 -1375 46
rect -1409 -46 -1375 -30
rect -1313 30 -1279 46
rect -1313 -46 -1279 -30
rect -1217 30 -1183 46
rect -1217 -46 -1183 -30
rect -1121 30 -1087 46
rect -1121 -46 -1087 -30
rect -1025 30 -991 46
rect -1025 -46 -991 -30
rect -929 30 -895 46
rect -929 -46 -895 -30
rect -833 30 -799 46
rect -833 -46 -799 -30
rect -737 30 -703 46
rect -737 -46 -703 -30
rect -641 30 -607 46
rect -641 -46 -607 -30
rect -545 30 -511 46
rect -545 -46 -511 -30
rect -449 30 -415 46
rect -449 -46 -415 -30
rect -353 30 -319 46
rect -353 -46 -319 -30
rect -257 30 -223 46
rect -257 -46 -223 -30
rect -161 30 -127 46
rect -161 -46 -127 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 127 30 161 46
rect 127 -46 161 -30
rect 223 30 257 46
rect 223 -46 257 -30
rect 319 30 353 46
rect 319 -46 353 -30
rect 415 30 449 46
rect 415 -46 449 -30
rect 511 30 545 46
rect 511 -46 545 -30
rect 607 30 641 46
rect 607 -46 641 -30
rect 703 30 737 46
rect 703 -46 737 -30
rect 799 30 833 46
rect 799 -46 833 -30
rect 895 30 929 46
rect 895 -46 929 -30
rect 991 30 1025 46
rect 991 -46 1025 -30
rect 1087 30 1121 46
rect 1087 -46 1121 -30
rect 1183 30 1217 46
rect 1183 -46 1217 -30
rect 1279 30 1313 46
rect 1279 -46 1313 -30
rect 1375 30 1409 46
rect 1375 -46 1409 -30
rect 1471 30 1505 46
rect 1471 -46 1505 -30
rect 1567 30 1601 46
rect 1567 -46 1601 -30
rect 1663 30 1697 46
rect 1663 -46 1697 -30
rect -1665 -123 -1649 -89
rect -1615 -123 -1599 -89
rect -1473 -123 -1457 -89
rect -1423 -123 -1407 -89
rect -1281 -123 -1265 -89
rect -1231 -123 -1215 -89
rect -1089 -123 -1073 -89
rect -1039 -123 -1023 -89
rect -897 -123 -881 -89
rect -847 -123 -831 -89
rect -705 -123 -689 -89
rect -655 -123 -639 -89
rect -513 -123 -497 -89
rect -463 -123 -447 -89
rect -321 -123 -305 -89
rect -271 -123 -255 -89
rect -129 -123 -113 -89
rect -79 -123 -63 -89
rect 63 -123 79 -89
rect 113 -123 129 -89
rect 255 -123 271 -89
rect 305 -123 321 -89
rect 447 -123 463 -89
rect 497 -123 513 -89
rect 639 -123 655 -89
rect 689 -123 705 -89
rect 831 -123 847 -89
rect 881 -123 897 -89
rect 1023 -123 1039 -89
rect 1073 -123 1089 -89
rect 1215 -123 1231 -89
rect 1265 -123 1281 -89
rect 1407 -123 1423 -89
rect 1457 -123 1473 -89
rect 1599 -123 1615 -89
rect 1649 -123 1665 -89
<< viali >>
rect -1697 -30 -1663 30
rect -1601 -30 -1567 30
rect -1505 -30 -1471 30
rect -1409 -30 -1375 30
rect -1313 -30 -1279 30
rect -1217 -30 -1183 30
rect -1121 -30 -1087 30
rect -1025 -30 -991 30
rect -929 -30 -895 30
rect -833 -30 -799 30
rect -737 -30 -703 30
rect -641 -30 -607 30
rect -545 -30 -511 30
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
rect 511 -30 545 30
rect 607 -30 641 30
rect 703 -30 737 30
rect 799 -30 833 30
rect 895 -30 929 30
rect 991 -30 1025 30
rect 1087 -30 1121 30
rect 1183 -30 1217 30
rect 1279 -30 1313 30
rect 1375 -30 1409 30
rect 1471 -30 1505 30
rect 1567 -30 1601 30
rect 1663 -30 1697 30
<< metal1 >>
rect -1703 30 -1657 42
rect -1703 -30 -1697 30
rect -1663 -30 -1657 30
rect -1703 -42 -1657 -30
rect -1607 30 -1561 42
rect -1607 -30 -1601 30
rect -1567 -30 -1561 30
rect -1607 -42 -1561 -30
rect -1511 30 -1465 42
rect -1511 -30 -1505 30
rect -1471 -30 -1465 30
rect -1511 -42 -1465 -30
rect -1415 30 -1369 42
rect -1415 -30 -1409 30
rect -1375 -30 -1369 30
rect -1415 -42 -1369 -30
rect -1319 30 -1273 42
rect -1319 -30 -1313 30
rect -1279 -30 -1273 30
rect -1319 -42 -1273 -30
rect -1223 30 -1177 42
rect -1223 -30 -1217 30
rect -1183 -30 -1177 30
rect -1223 -42 -1177 -30
rect -1127 30 -1081 42
rect -1127 -30 -1121 30
rect -1087 -30 -1081 30
rect -1127 -42 -1081 -30
rect -1031 30 -985 42
rect -1031 -30 -1025 30
rect -991 -30 -985 30
rect -1031 -42 -985 -30
rect -935 30 -889 42
rect -935 -30 -929 30
rect -895 -30 -889 30
rect -935 -42 -889 -30
rect -839 30 -793 42
rect -839 -30 -833 30
rect -799 -30 -793 30
rect -839 -42 -793 -30
rect -743 30 -697 42
rect -743 -30 -737 30
rect -703 -30 -697 30
rect -743 -42 -697 -30
rect -647 30 -601 42
rect -647 -30 -641 30
rect -607 -30 -601 30
rect -647 -42 -601 -30
rect -551 30 -505 42
rect -551 -30 -545 30
rect -511 -30 -505 30
rect -551 -42 -505 -30
rect -455 30 -409 42
rect -455 -30 -449 30
rect -415 -30 -409 30
rect -455 -42 -409 -30
rect -359 30 -313 42
rect -359 -30 -353 30
rect -319 -30 -313 30
rect -359 -42 -313 -30
rect -263 30 -217 42
rect -263 -30 -257 30
rect -223 -30 -217 30
rect -263 -42 -217 -30
rect -167 30 -121 42
rect -167 -30 -161 30
rect -127 -30 -121 30
rect -167 -42 -121 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 121 30 167 42
rect 121 -30 127 30
rect 161 -30 167 30
rect 121 -42 167 -30
rect 217 30 263 42
rect 217 -30 223 30
rect 257 -30 263 30
rect 217 -42 263 -30
rect 313 30 359 42
rect 313 -30 319 30
rect 353 -30 359 30
rect 313 -42 359 -30
rect 409 30 455 42
rect 409 -30 415 30
rect 449 -30 455 30
rect 409 -42 455 -30
rect 505 30 551 42
rect 505 -30 511 30
rect 545 -30 551 30
rect 505 -42 551 -30
rect 601 30 647 42
rect 601 -30 607 30
rect 641 -30 647 30
rect 601 -42 647 -30
rect 697 30 743 42
rect 697 -30 703 30
rect 737 -30 743 30
rect 697 -42 743 -30
rect 793 30 839 42
rect 793 -30 799 30
rect 833 -30 839 30
rect 793 -42 839 -30
rect 889 30 935 42
rect 889 -30 895 30
rect 929 -30 935 30
rect 889 -42 935 -30
rect 985 30 1031 42
rect 985 -30 991 30
rect 1025 -30 1031 30
rect 985 -42 1031 -30
rect 1081 30 1127 42
rect 1081 -30 1087 30
rect 1121 -30 1127 30
rect 1081 -42 1127 -30
rect 1177 30 1223 42
rect 1177 -30 1183 30
rect 1217 -30 1223 30
rect 1177 -42 1223 -30
rect 1273 30 1319 42
rect 1273 -30 1279 30
rect 1313 -30 1319 30
rect 1273 -42 1319 -30
rect 1369 30 1415 42
rect 1369 -30 1375 30
rect 1409 -30 1415 30
rect 1369 -42 1415 -30
rect 1465 30 1511 42
rect 1465 -30 1471 30
rect 1505 -30 1511 30
rect 1465 -42 1511 -30
rect 1561 30 1607 42
rect 1561 -30 1567 30
rect 1601 -30 1607 30
rect 1561 -42 1607 -30
rect 1657 30 1703 42
rect 1657 -30 1663 30
rect 1697 -30 1703 30
rect 1657 -42 1703 -30
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 35 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
