magic
tech sky130A
magscale 1 2
timestamp 1698179620
<< error_s >>
rect -1230 3631 -1088 3652
rect -1202 3603 -1116 3624
<< locali >>
rect 488 4848 562 4932
rect 474 3738 562 3830
rect 474 3730 600 3738
rect -1406 3234 -1347 3381
rect -2215 2557 -1907 2591
rect -1827 2545 -1682 2579
rect -1440 2562 -1295 2596
rect -1059 2549 -751 2583
rect -2032 2386 -1991 2491
rect -867 2386 -826 2491
rect -2255 2365 -599 2386
rect -2255 2308 -599 2325
<< viali >>
rect -2255 2325 -599 2365
<< metal1 >>
rect -3151 4838 -2789 4873
rect -3151 3456 -3116 4838
rect 54 4678 64 4744
rect 152 4678 162 4744
rect 3506 4678 3516 4738
rect 3622 4678 3632 4738
rect -1190 4552 -1180 4632
rect -1102 4552 -1092 4632
rect -3042 3945 -2810 3986
rect -3042 3580 -3001 3945
rect -1922 3604 -1912 3666
rect -1836 3604 -1826 3666
rect 736 3620 746 3676
rect 830 3620 840 3676
rect -3042 3539 -1955 3580
rect -3151 3421 -2232 3456
rect -2267 2386 -2232 3421
rect -1996 2904 -1955 3539
rect -1914 2998 -1877 3604
rect -1212 3516 -1202 3614
rect -1116 3516 -1106 3614
rect -1212 3129 -1175 3516
rect -1808 3061 -1254 3098
rect -1914 2990 -1112 2998
rect -1914 2961 1286 2990
rect -1149 2958 1286 2961
rect -1996 2863 -1541 2904
rect -1551 2822 -1541 2863
rect -1452 2822 -1442 2904
rect -1712 2672 -1702 2740
rect -1594 2672 -1584 2740
rect -1542 2544 -1501 2822
rect -1149 2542 -1112 2958
rect -630 2802 -620 2892
rect -530 2802 -520 2892
rect 1254 2662 1286 2958
rect 1254 2630 1874 2662
rect 1842 2532 1874 2630
rect 2162 2530 2172 2584
rect 2238 2530 2248 2584
rect -1683 2433 -1673 2495
rect -1566 2481 -1556 2495
rect -1566 2452 -1201 2481
rect -1566 2433 -1556 2452
rect -2267 2371 -599 2386
rect -2267 2365 -587 2371
rect -2267 2325 -2255 2365
rect -599 2353 -587 2365
rect -599 2325 -143 2353
rect -2432 2259 -2422 2320
rect -2362 2259 -2352 2320
rect -2267 2319 -143 2325
rect -2255 2316 -143 2319
rect -2255 2308 -599 2316
rect -180 1883 -143 2316
rect -203 1824 -193 1883
rect -130 1824 -120 1883
<< via1 >>
rect 64 4678 152 4744
rect 3516 4678 3622 4738
rect -1180 4552 -1102 4632
rect -1912 3604 -1836 3666
rect 746 3620 830 3676
rect -1202 3516 -1116 3614
rect -1541 2822 -1452 2904
rect -1702 2672 -1594 2740
rect -620 2802 -530 2892
rect 2172 2530 2238 2584
rect -1673 2433 -1566 2495
rect -2422 2259 -2362 2320
rect -193 1824 -130 1883
<< metal2 >>
rect -3283 5005 -1134 5043
rect -3283 2764 -3245 5005
rect -1172 4642 -1134 5005
rect 68 4998 3572 5054
rect 68 4754 124 4998
rect 64 4744 152 4754
rect 64 4668 152 4678
rect 3516 4748 3572 4998
rect 3516 4738 3622 4748
rect 3516 4668 3622 4678
rect -1180 4632 -1102 4642
rect -1180 4542 -1102 4552
rect -2189 3672 -2147 4199
rect 746 3681 830 3686
rect 491 3676 830 3681
rect -1912 3672 -1836 3676
rect -2192 3666 -1836 3672
rect -2192 3630 -1912 3666
rect 491 3639 746 3676
rect -1912 3594 -1836 3604
rect -1202 3614 -1116 3624
rect -1208 3526 -1202 3568
rect 491 3568 533 3639
rect 746 3610 830 3620
rect -1116 3526 533 3568
rect -1202 3506 -1116 3516
rect 1116 3382 1144 4054
rect -1541 2904 -1452 2914
rect -620 2892 -530 2902
rect -1452 2822 -620 2876
rect -1541 2812 -1452 2822
rect -620 2792 -530 2802
rect -3283 2750 -1614 2764
rect -3283 2740 -1594 2750
rect -3283 2728 -1702 2740
rect -3283 2727 -3245 2728
rect -1702 2662 -1594 2672
rect 2172 2588 2238 2598
rect 2172 2520 2238 2530
rect -1673 2495 -1566 2505
rect -2367 2442 -1673 2481
rect -2367 2341 -2328 2442
rect -1673 2423 -1566 2433
rect -2442 2331 -2328 2341
rect -2340 2285 -2328 2331
rect -2442 2232 -2340 2242
rect -213 1890 -129 1900
rect -213 1796 -129 1806
<< via2 >>
rect -620 2802 -530 2892
rect 2172 2584 2238 2588
rect 2172 2530 2238 2584
rect -2442 2320 -2340 2331
rect -2442 2259 -2422 2320
rect -2422 2259 -2362 2320
rect -2362 2259 -2340 2320
rect -2442 2242 -2340 2259
rect -213 1883 -129 1890
rect -213 1824 -193 1883
rect -193 1824 -130 1883
rect -130 1824 -129 1883
rect -213 1806 -129 1824
<< metal3 >>
rect -630 2892 -520 2897
rect -630 2802 -620 2892
rect -530 2866 -520 2892
rect -530 2806 2266 2866
rect -530 2802 -520 2806
rect -630 2797 -520 2802
rect 2206 2593 2266 2806
rect 2162 2588 2266 2593
rect 2162 2530 2172 2588
rect 2238 2530 2266 2588
rect 2162 2525 2248 2530
rect -2474 2214 -2464 2376
rect -2314 2214 -2304 2376
rect -223 1890 -119 1895
rect -223 1806 -213 1890
rect -129 1806 -119 1890
rect -223 1801 -119 1806
<< via3 >>
rect -2464 2331 -2314 2376
rect -2464 2242 -2442 2331
rect -2442 2242 -2340 2331
rect -2340 2242 -2314 2331
rect -2464 2214 -2314 2242
<< metal4 >>
rect -2465 2376 -2313 2377
rect -2465 2214 -2464 2376
rect -2314 2273 -2313 2376
rect -2314 2214 -2300 2273
rect -2465 2213 -2300 2214
rect -2363 1940 -2300 2213
use cmfb  cmfb_0
timestamp 1698179620
transform 1 0 -3134 0 1 2875
box 203 439 3639 2056
use integrator_full_new1  integrator_full_new1_0
timestamp 1698179620
transform 1 0 386 0 1 3314
box -386 -3314 3986 1624
use sky130_fd_pr__nfet_01v8_53744R  sky130_fd_pr__nfet_01v8_53744R_0
timestamp 1698166690
transform 0 1 -1344 -1 0 3174
box -246 -310 246 310
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_0
timestamp 1698155087
transform 1 0 -1233 0 1 2582
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_1
timestamp 1698155087
transform 1 0 -1619 0 1 2582
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_2
timestamp 1698155087
transform 1 0 -2005 0 1 2582
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_3
timestamp 1698155087
transform 1 0 -847 0 1 2582
box -246 -269 246 269
use sky130_fd_pr__cap_mim_m3_1_4PHTN9  XC3
timestamp 1697610037
transform 1 0 -1291 0 1 1094
box -1186 -1040 1186 1040
<< end >>
