magic
tech sky130A
magscale 1 2
timestamp 1697695294
<< error_p >>
rect -29 114 29 120
rect -29 80 -17 114
rect -29 74 29 80
rect -125 -80 -67 -74
rect 67 -80 125 -74
rect -125 -114 -113 -80
rect 67 -114 79 -80
rect -125 -120 -67 -114
rect 67 -120 125 -114
<< nmos >>
rect -111 -42 -81 42
rect -15 -42 15 42
rect 81 -42 111 42
<< ndiff >>
rect -173 30 -111 42
rect -173 -30 -161 30
rect -127 -30 -111 30
rect -173 -42 -111 -30
rect -81 30 -15 42
rect -81 -30 -65 30
rect -31 -30 -15 30
rect -81 -42 -15 -30
rect 15 30 81 42
rect 15 -30 31 30
rect 65 -30 81 30
rect 15 -42 81 -30
rect 111 30 173 42
rect 111 -30 127 30
rect 161 -30 173 30
rect 111 -42 173 -30
<< ndiffc >>
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
<< poly >>
rect -33 114 33 130
rect -33 80 -17 114
rect 17 80 33 114
rect -111 42 -81 68
rect -33 64 33 80
rect -15 42 15 64
rect 81 42 111 68
rect -111 -64 -81 -42
rect -129 -80 -63 -64
rect -15 -68 15 -42
rect 81 -64 111 -42
rect -129 -114 -113 -80
rect -79 -114 -63 -80
rect -129 -130 -63 -114
rect 63 -80 129 -64
rect 63 -114 79 -80
rect 113 -114 129 -80
rect 63 -130 129 -114
<< polycont >>
rect -17 80 17 114
rect -113 -114 -79 -80
rect 79 -114 113 -80
<< locali >>
rect -33 80 -17 114
rect 17 80 33 114
rect -161 30 -127 46
rect -161 -46 -127 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 127 30 161 46
rect 127 -46 161 -30
rect -129 -114 -113 -80
rect -79 -114 -63 -80
rect 63 -114 79 -80
rect 113 -114 129 -80
<< viali >>
rect -17 80 17 114
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect -113 -114 -79 -80
rect 79 -114 113 -80
<< metal1 >>
rect -29 114 29 120
rect -29 80 -17 114
rect 17 80 29 114
rect -29 74 29 80
rect -167 30 -121 42
rect -167 -30 -161 30
rect -127 -30 -121 30
rect -167 -42 -121 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 121 30 167 42
rect 121 -30 127 30
rect 161 -30 167 30
rect 121 -42 167 -30
rect -125 -80 -67 -74
rect -125 -114 -113 -80
rect -79 -114 -67 -80
rect -125 -120 -67 -114
rect 67 -80 125 -74
rect 67 -114 79 -80
rect 113 -114 125 -80
rect 67 -120 125 -114
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
