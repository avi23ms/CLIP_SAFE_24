magic
tech sky130A
magscale 1 2
timestamp 1699103691
<< nmos >>
rect -1263 -42 -1233 42
rect -1167 -42 -1137 42
rect -1071 -42 -1041 42
rect -975 -42 -945 42
rect -879 -42 -849 42
rect -783 -42 -753 42
rect -687 -42 -657 42
rect -591 -42 -561 42
rect -495 -42 -465 42
rect -399 -42 -369 42
rect -303 -42 -273 42
rect -207 -42 -177 42
rect -111 -42 -81 42
rect -15 -42 15 42
rect 81 -42 111 42
rect 177 -42 207 42
rect 273 -42 303 42
rect 369 -42 399 42
rect 465 -42 495 42
rect 561 -42 591 42
rect 657 -42 687 42
rect 753 -42 783 42
rect 849 -42 879 42
rect 945 -42 975 42
rect 1041 -42 1071 42
rect 1137 -42 1167 42
rect 1233 -42 1263 42
<< ndiff >>
rect -1325 30 -1263 42
rect -1325 -30 -1313 30
rect -1279 -30 -1263 30
rect -1325 -42 -1263 -30
rect -1233 30 -1167 42
rect -1233 -30 -1217 30
rect -1183 -30 -1167 30
rect -1233 -42 -1167 -30
rect -1137 30 -1071 42
rect -1137 -30 -1121 30
rect -1087 -30 -1071 30
rect -1137 -42 -1071 -30
rect -1041 30 -975 42
rect -1041 -30 -1025 30
rect -991 -30 -975 30
rect -1041 -42 -975 -30
rect -945 30 -879 42
rect -945 -30 -929 30
rect -895 -30 -879 30
rect -945 -42 -879 -30
rect -849 30 -783 42
rect -849 -30 -833 30
rect -799 -30 -783 30
rect -849 -42 -783 -30
rect -753 30 -687 42
rect -753 -30 -737 30
rect -703 -30 -687 30
rect -753 -42 -687 -30
rect -657 30 -591 42
rect -657 -30 -641 30
rect -607 -30 -591 30
rect -657 -42 -591 -30
rect -561 30 -495 42
rect -561 -30 -545 30
rect -511 -30 -495 30
rect -561 -42 -495 -30
rect -465 30 -399 42
rect -465 -30 -449 30
rect -415 -30 -399 30
rect -465 -42 -399 -30
rect -369 30 -303 42
rect -369 -30 -353 30
rect -319 -30 -303 30
rect -369 -42 -303 -30
rect -273 30 -207 42
rect -273 -30 -257 30
rect -223 -30 -207 30
rect -273 -42 -207 -30
rect -177 30 -111 42
rect -177 -30 -161 30
rect -127 -30 -111 30
rect -177 -42 -111 -30
rect -81 30 -15 42
rect -81 -30 -65 30
rect -31 -30 -15 30
rect -81 -42 -15 -30
rect 15 30 81 42
rect 15 -30 31 30
rect 65 -30 81 30
rect 15 -42 81 -30
rect 111 30 177 42
rect 111 -30 127 30
rect 161 -30 177 30
rect 111 -42 177 -30
rect 207 30 273 42
rect 207 -30 223 30
rect 257 -30 273 30
rect 207 -42 273 -30
rect 303 30 369 42
rect 303 -30 319 30
rect 353 -30 369 30
rect 303 -42 369 -30
rect 399 30 465 42
rect 399 -30 415 30
rect 449 -30 465 30
rect 399 -42 465 -30
rect 495 30 561 42
rect 495 -30 511 30
rect 545 -30 561 30
rect 495 -42 561 -30
rect 591 30 657 42
rect 591 -30 607 30
rect 641 -30 657 30
rect 591 -42 657 -30
rect 687 30 753 42
rect 687 -30 703 30
rect 737 -30 753 30
rect 687 -42 753 -30
rect 783 30 849 42
rect 783 -30 799 30
rect 833 -30 849 30
rect 783 -42 849 -30
rect 879 30 945 42
rect 879 -30 895 30
rect 929 -30 945 30
rect 879 -42 945 -30
rect 975 30 1041 42
rect 975 -30 991 30
rect 1025 -30 1041 30
rect 975 -42 1041 -30
rect 1071 30 1137 42
rect 1071 -30 1087 30
rect 1121 -30 1137 30
rect 1071 -42 1137 -30
rect 1167 30 1233 42
rect 1167 -30 1183 30
rect 1217 -30 1233 30
rect 1167 -42 1233 -30
rect 1263 30 1325 42
rect 1263 -30 1279 30
rect 1313 -30 1325 30
rect 1263 -42 1325 -30
<< ndiffc >>
rect -1313 -30 -1279 30
rect -1217 -30 -1183 30
rect -1121 -30 -1087 30
rect -1025 -30 -991 30
rect -929 -30 -895 30
rect -833 -30 -799 30
rect -737 -30 -703 30
rect -641 -30 -607 30
rect -545 -30 -511 30
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
rect 511 -30 545 30
rect 607 -30 641 30
rect 703 -30 737 30
rect 799 -30 833 30
rect 895 -30 929 30
rect 991 -30 1025 30
rect 1087 -30 1121 30
rect 1183 -30 1217 30
rect 1279 -30 1313 30
<< poly >>
rect -1185 114 -1119 130
rect -1185 80 -1169 114
rect -1135 80 -1119 114
rect -1263 42 -1233 68
rect -1185 64 -1119 80
rect -993 114 -927 130
rect -993 80 -977 114
rect -943 80 -927 114
rect -1167 42 -1137 64
rect -1071 42 -1041 68
rect -993 64 -927 80
rect -801 114 -735 130
rect -801 80 -785 114
rect -751 80 -735 114
rect -975 42 -945 64
rect -879 42 -849 68
rect -801 64 -735 80
rect -609 114 -543 130
rect -609 80 -593 114
rect -559 80 -543 114
rect -783 42 -753 64
rect -687 42 -657 68
rect -609 64 -543 80
rect -417 114 -351 130
rect -417 80 -401 114
rect -367 80 -351 114
rect -591 42 -561 64
rect -495 42 -465 68
rect -417 64 -351 80
rect -225 114 -159 130
rect -225 80 -209 114
rect -175 80 -159 114
rect -399 42 -369 64
rect -303 42 -273 68
rect -225 64 -159 80
rect -33 114 33 130
rect -33 80 -17 114
rect 17 80 33 114
rect -207 42 -177 64
rect -111 42 -81 68
rect -33 64 33 80
rect 159 114 225 130
rect 159 80 175 114
rect 209 80 225 114
rect -15 42 15 64
rect 81 42 111 68
rect 159 64 225 80
rect 351 114 417 130
rect 351 80 367 114
rect 401 80 417 114
rect 177 42 207 64
rect 273 42 303 68
rect 351 64 417 80
rect 543 114 609 130
rect 543 80 559 114
rect 593 80 609 114
rect 369 42 399 64
rect 465 42 495 68
rect 543 64 609 80
rect 735 114 801 130
rect 735 80 751 114
rect 785 80 801 114
rect 561 42 591 64
rect 657 42 687 68
rect 735 64 801 80
rect 927 114 993 130
rect 927 80 943 114
rect 977 80 993 114
rect 753 42 783 64
rect 849 42 879 68
rect 927 64 993 80
rect 1119 114 1185 130
rect 1119 80 1135 114
rect 1169 80 1185 114
rect 945 42 975 64
rect 1041 42 1071 68
rect 1119 64 1185 80
rect 1137 42 1167 64
rect 1233 42 1263 68
rect -1263 -64 -1233 -42
rect -1281 -80 -1215 -64
rect -1167 -68 -1137 -42
rect -1071 -64 -1041 -42
rect -1281 -114 -1265 -80
rect -1231 -114 -1215 -80
rect -1281 -130 -1215 -114
rect -1089 -80 -1023 -64
rect -975 -68 -945 -42
rect -879 -64 -849 -42
rect -1089 -114 -1073 -80
rect -1039 -114 -1023 -80
rect -1089 -130 -1023 -114
rect -897 -80 -831 -64
rect -783 -68 -753 -42
rect -687 -64 -657 -42
rect -897 -114 -881 -80
rect -847 -114 -831 -80
rect -897 -130 -831 -114
rect -705 -80 -639 -64
rect -591 -68 -561 -42
rect -495 -64 -465 -42
rect -705 -114 -689 -80
rect -655 -114 -639 -80
rect -705 -130 -639 -114
rect -513 -80 -447 -64
rect -399 -68 -369 -42
rect -303 -64 -273 -42
rect -513 -114 -497 -80
rect -463 -114 -447 -80
rect -513 -130 -447 -114
rect -321 -80 -255 -64
rect -207 -68 -177 -42
rect -111 -64 -81 -42
rect -321 -114 -305 -80
rect -271 -114 -255 -80
rect -321 -130 -255 -114
rect -129 -80 -63 -64
rect -15 -68 15 -42
rect 81 -64 111 -42
rect -129 -114 -113 -80
rect -79 -114 -63 -80
rect -129 -130 -63 -114
rect 63 -80 129 -64
rect 177 -68 207 -42
rect 273 -64 303 -42
rect 63 -114 79 -80
rect 113 -114 129 -80
rect 63 -130 129 -114
rect 255 -80 321 -64
rect 369 -68 399 -42
rect 465 -64 495 -42
rect 255 -114 271 -80
rect 305 -114 321 -80
rect 255 -130 321 -114
rect 447 -80 513 -64
rect 561 -68 591 -42
rect 657 -64 687 -42
rect 447 -114 463 -80
rect 497 -114 513 -80
rect 447 -130 513 -114
rect 639 -80 705 -64
rect 753 -68 783 -42
rect 849 -64 879 -42
rect 639 -114 655 -80
rect 689 -114 705 -80
rect 639 -130 705 -114
rect 831 -80 897 -64
rect 945 -68 975 -42
rect 1041 -64 1071 -42
rect 831 -114 847 -80
rect 881 -114 897 -80
rect 831 -130 897 -114
rect 1023 -80 1089 -64
rect 1137 -68 1167 -42
rect 1233 -64 1263 -42
rect 1023 -114 1039 -80
rect 1073 -114 1089 -80
rect 1023 -130 1089 -114
rect 1215 -80 1281 -64
rect 1215 -114 1231 -80
rect 1265 -114 1281 -80
rect 1215 -130 1281 -114
<< polycont >>
rect -1169 80 -1135 114
rect -977 80 -943 114
rect -785 80 -751 114
rect -593 80 -559 114
rect -401 80 -367 114
rect -209 80 -175 114
rect -17 80 17 114
rect 175 80 209 114
rect 367 80 401 114
rect 559 80 593 114
rect 751 80 785 114
rect 943 80 977 114
rect 1135 80 1169 114
rect -1265 -114 -1231 -80
rect -1073 -114 -1039 -80
rect -881 -114 -847 -80
rect -689 -114 -655 -80
rect -497 -114 -463 -80
rect -305 -114 -271 -80
rect -113 -114 -79 -80
rect 79 -114 113 -80
rect 271 -114 305 -80
rect 463 -114 497 -80
rect 655 -114 689 -80
rect 847 -114 881 -80
rect 1039 -114 1073 -80
rect 1231 -114 1265 -80
<< locali >>
rect -1185 80 -1169 114
rect -1135 80 -1119 114
rect -993 80 -977 114
rect -943 80 -927 114
rect -801 80 -785 114
rect -751 80 -735 114
rect -609 80 -593 114
rect -559 80 -543 114
rect -417 80 -401 114
rect -367 80 -351 114
rect -225 80 -209 114
rect -175 80 -159 114
rect -33 80 -17 114
rect 17 80 33 114
rect 159 80 175 114
rect 209 80 225 114
rect 351 80 367 114
rect 401 80 417 114
rect 543 80 559 114
rect 593 80 609 114
rect 735 80 751 114
rect 785 80 801 114
rect 927 80 943 114
rect 977 80 993 114
rect 1119 80 1135 114
rect 1169 80 1185 114
rect -1313 30 -1279 46
rect -1313 -46 -1279 -30
rect -1217 30 -1183 46
rect -1217 -46 -1183 -30
rect -1121 30 -1087 46
rect -1121 -46 -1087 -30
rect -1025 30 -991 46
rect -1025 -46 -991 -30
rect -929 30 -895 46
rect -929 -46 -895 -30
rect -833 30 -799 46
rect -833 -46 -799 -30
rect -737 30 -703 46
rect -737 -46 -703 -30
rect -641 30 -607 46
rect -641 -46 -607 -30
rect -545 30 -511 46
rect -545 -46 -511 -30
rect -449 30 -415 46
rect -449 -46 -415 -30
rect -353 30 -319 46
rect -353 -46 -319 -30
rect -257 30 -223 46
rect -257 -46 -223 -30
rect -161 30 -127 46
rect -161 -46 -127 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 127 30 161 46
rect 127 -46 161 -30
rect 223 30 257 46
rect 223 -46 257 -30
rect 319 30 353 46
rect 319 -46 353 -30
rect 415 30 449 46
rect 415 -46 449 -30
rect 511 30 545 46
rect 511 -46 545 -30
rect 607 30 641 46
rect 607 -46 641 -30
rect 703 30 737 46
rect 703 -46 737 -30
rect 799 30 833 46
rect 799 -46 833 -30
rect 895 30 929 46
rect 895 -46 929 -30
rect 991 30 1025 46
rect 991 -46 1025 -30
rect 1087 30 1121 46
rect 1087 -46 1121 -30
rect 1183 30 1217 46
rect 1183 -46 1217 -30
rect 1279 30 1313 46
rect 1279 -46 1313 -30
rect -1281 -114 -1265 -80
rect -1231 -114 -1215 -80
rect -1089 -114 -1073 -80
rect -1039 -114 -1023 -80
rect -897 -114 -881 -80
rect -847 -114 -831 -80
rect -705 -114 -689 -80
rect -655 -114 -639 -80
rect -513 -114 -497 -80
rect -463 -114 -447 -80
rect -321 -114 -305 -80
rect -271 -114 -255 -80
rect -129 -114 -113 -80
rect -79 -114 -63 -80
rect 63 -114 79 -80
rect 113 -114 129 -80
rect 255 -114 271 -80
rect 305 -114 321 -80
rect 447 -114 463 -80
rect 497 -114 513 -80
rect 639 -114 655 -80
rect 689 -114 705 -80
rect 831 -114 847 -80
rect 881 -114 897 -80
rect 1023 -114 1039 -80
rect 1073 -114 1089 -80
rect 1215 -114 1231 -80
rect 1265 -114 1281 -80
<< viali >>
rect -1313 -30 -1279 30
rect -1217 -30 -1183 30
rect -1121 -30 -1087 30
rect -1025 -30 -991 30
rect -929 -30 -895 30
rect -833 -30 -799 30
rect -737 -30 -703 30
rect -641 -30 -607 30
rect -545 -30 -511 30
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
rect 511 -30 545 30
rect 607 -30 641 30
rect 703 -30 737 30
rect 799 -30 833 30
rect 895 -30 929 30
rect 991 -30 1025 30
rect 1087 -30 1121 30
rect 1183 -30 1217 30
rect 1279 -30 1313 30
<< metal1 >>
rect -1319 30 -1273 42
rect -1319 -30 -1313 30
rect -1279 -30 -1273 30
rect -1319 -42 -1273 -30
rect -1223 30 -1177 42
rect -1223 -30 -1217 30
rect -1183 -30 -1177 30
rect -1223 -42 -1177 -30
rect -1127 30 -1081 42
rect -1127 -30 -1121 30
rect -1087 -30 -1081 30
rect -1127 -42 -1081 -30
rect -1031 30 -985 42
rect -1031 -30 -1025 30
rect -991 -30 -985 30
rect -1031 -42 -985 -30
rect -935 30 -889 42
rect -935 -30 -929 30
rect -895 -30 -889 30
rect -935 -42 -889 -30
rect -839 30 -793 42
rect -839 -30 -833 30
rect -799 -30 -793 30
rect -839 -42 -793 -30
rect -743 30 -697 42
rect -743 -30 -737 30
rect -703 -30 -697 30
rect -743 -42 -697 -30
rect -647 30 -601 42
rect -647 -30 -641 30
rect -607 -30 -601 30
rect -647 -42 -601 -30
rect -551 30 -505 42
rect -551 -30 -545 30
rect -511 -30 -505 30
rect -551 -42 -505 -30
rect -455 30 -409 42
rect -455 -30 -449 30
rect -415 -30 -409 30
rect -455 -42 -409 -30
rect -359 30 -313 42
rect -359 -30 -353 30
rect -319 -30 -313 30
rect -359 -42 -313 -30
rect -263 30 -217 42
rect -263 -30 -257 30
rect -223 -30 -217 30
rect -263 -42 -217 -30
rect -167 30 -121 42
rect -167 -30 -161 30
rect -127 -30 -121 30
rect -167 -42 -121 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 121 30 167 42
rect 121 -30 127 30
rect 161 -30 167 30
rect 121 -42 167 -30
rect 217 30 263 42
rect 217 -30 223 30
rect 257 -30 263 30
rect 217 -42 263 -30
rect 313 30 359 42
rect 313 -30 319 30
rect 353 -30 359 30
rect 313 -42 359 -30
rect 409 30 455 42
rect 409 -30 415 30
rect 449 -30 455 30
rect 409 -42 455 -30
rect 505 30 551 42
rect 505 -30 511 30
rect 545 -30 551 30
rect 505 -42 551 -30
rect 601 30 647 42
rect 601 -30 607 30
rect 641 -30 647 30
rect 601 -42 647 -30
rect 697 30 743 42
rect 697 -30 703 30
rect 737 -30 743 30
rect 697 -42 743 -30
rect 793 30 839 42
rect 793 -30 799 30
rect 833 -30 839 30
rect 793 -42 839 -30
rect 889 30 935 42
rect 889 -30 895 30
rect 929 -30 935 30
rect 889 -42 935 -30
rect 985 30 1031 42
rect 985 -30 991 30
rect 1025 -30 1031 30
rect 985 -42 1031 -30
rect 1081 30 1127 42
rect 1081 -30 1087 30
rect 1121 -30 1127 30
rect 1081 -42 1127 -30
rect 1177 30 1223 42
rect 1177 -30 1183 30
rect 1217 -30 1223 30
rect 1177 -42 1223 -30
rect 1273 30 1319 42
rect 1273 -30 1279 30
rect 1313 -30 1319 30
rect 1273 -42 1319 -30
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 27 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
