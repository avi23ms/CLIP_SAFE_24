magic
tech sky130A
magscale 1 2
timestamp 1698684236
<< error_s >>
rect 16120 14494 16711 14496
rect 15906 14492 16711 14494
rect 15615 14488 16711 14492
rect 16096 12408 16703 12410
rect 15882 12406 16703 12408
rect 15607 12404 16703 12406
rect 8361 12400 8948 12402
rect 8361 12398 9162 12400
rect 8361 12394 9457 12398
rect 8365 10314 8940 10316
rect 8365 10312 9154 10314
rect 8365 10310 9461 10312
rect 8357 8228 8930 8230
rect 8357 8226 9144 8228
rect 8357 8224 9453 8226
rect 16112 8208 16735 8210
rect 8347 6142 8930 6144
rect 8347 6140 9144 6142
rect 8347 6138 9443 6140
rect 16048 6124 16695 6126
rect 15834 6122 16695 6124
rect 15599 6118 16695 6122
rect 8347 4058 8942 4060
rect 8347 4056 9156 4058
rect 8347 4052 9443 4056
rect 16026 4038 16631 4040
rect 15812 4036 16631 4038
rect 15535 4034 16631 4036
rect 2526 2326 2570 2340
rect 2710 2338 2760 2340
rect 2806 2338 2856 2340
rect 2902 2338 2952 2340
rect 2998 2338 3048 2340
rect 3094 2338 3144 2340
rect 3190 2338 3240 2340
rect 3286 2338 3336 2340
rect 3382 2338 3432 2340
rect 3478 2338 3528 2340
rect 3574 2338 3624 2340
rect 3670 2338 3720 2340
rect 3766 2338 3816 2340
rect 3862 2338 3912 2340
rect 3958 2338 4008 2340
rect 4054 2338 4104 2340
rect 4150 2338 4200 2340
rect 4246 2338 4296 2340
rect 4342 2338 4392 2340
rect 4438 2338 4488 2340
rect 4534 2338 4584 2340
rect 16029 1954 16609 1956
rect 15815 1952 16609 1954
rect 15513 1948 16609 1952
rect 15605 272 16499 274
rect 15577 244 16527 246
rect 15533 194 16595 202
rect 15503 186 16649 194
rect 16661 186 17749 192
rect 15561 166 15607 174
rect 15657 166 15703 174
rect 15753 166 15799 174
rect 15849 166 15895 174
rect 15945 166 15991 174
rect 16041 166 16087 174
rect 16137 166 16183 174
rect 16233 166 16279 174
rect 16329 166 16375 174
rect 16425 166 16471 174
rect 16521 166 16567 174
rect 15531 158 16621 166
rect 16689 158 17721 164
rect 20300 22 20341 38
rect 20328 -6 20341 10
<< psubdiff >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
<< nsubdiff >>
rect 12396 17402 12508 17434
rect 12396 17294 12430 17402
rect 12484 17294 12508 17402
rect 12396 17274 12508 17294
<< psubdiffcont >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
<< nsubdiffcont >>
rect 12430 17294 12484 17402
<< locali >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
rect 12396 17402 12506 17436
rect 12396 17294 12430 17402
rect 12484 17294 12506 17402
rect 12396 17262 12506 17294
<< viali >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 12430 17294 12484 17402
<< metal1 >>
rect 12288 19430 12324 19490
rect 13062 19440 13098 19554
rect 12200 19428 12324 19430
rect 1010 19426 12324 19428
rect 946 19396 12324 19426
rect 13052 19414 13220 19440
rect 23646 19414 24070 19418
rect 946 19260 12330 19396
rect 946 19238 12324 19260
rect 13052 19246 24070 19414
rect 13052 19240 13220 19246
rect 946 19235 12317 19238
rect 946 17770 1204 19235
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
rect 12370 18132 12534 18148
rect 946 17412 970 17770
rect 1172 17412 1204 17770
rect 946 17386 1204 17412
rect 12370 17290 12400 18132
rect 12502 17290 12534 18132
rect 23646 17930 24070 19246
rect 14430 17600 14534 17698
rect 14430 17508 14720 17600
rect 23646 17488 23674 17930
rect 24008 17488 24070 17930
rect 23646 17444 24070 17488
rect 12370 17240 12534 17290
rect 4517 254 12354 258
rect 4360 172 12354 254
rect 12660 188 20476 246
rect 12660 186 20478 188
rect 4360 32 4904 172
rect 19196 156 20478 186
rect 4360 -324 4412 32
rect 4854 -324 4904 32
rect 4360 -374 4904 -324
rect 12464 108 12550 120
rect 4541 -377 4627 -374
rect 12464 -472 12478 108
rect 12538 -472 12550 108
rect 19196 52 19222 156
rect 20440 52 20478 156
rect 19196 22 20478 52
rect 20410 -122 20470 22
rect 12464 -576 12550 -472
rect 936 -701 1482 -688
rect 8366 -701 8664 -698
rect 936 -735 8838 -701
rect 23632 -706 24074 -694
rect 936 -788 1482 -735
rect 936 -1984 1006 -788
rect 1406 -1984 1482 -788
rect 8366 -744 8664 -735
rect 16128 -742 24074 -706
rect 8366 -1102 8398 -744
rect 8632 -1102 8664 -744
rect 8366 -1446 8664 -1102
rect 16224 -750 16610 -742
rect 16224 -1082 16268 -750
rect 16572 -1082 16610 -750
rect 16224 -1464 16610 -1082
rect 23632 -752 24074 -742
rect 23632 -1826 23696 -752
rect 23998 -1826 24074 -752
rect 23632 -1902 24074 -1826
rect 936 -2064 1482 -1984
<< via1 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 970 17412 1172 17770
rect 12400 17402 12502 18132
rect 12400 17294 12430 17402
rect 12430 17294 12484 17402
rect 12484 17294 12502 17402
rect 12400 17290 12502 17294
rect 23674 17488 24008 17930
rect 4412 -324 4854 32
rect 12478 -472 12538 108
rect 19222 52 20440 156
rect 1006 -1984 1406 -788
rect 8398 -1102 8632 -744
rect 16268 -1082 16572 -750
rect 23696 -1826 23998 -752
<< metal2 >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
rect 12370 18132 12540 18174
rect 946 17770 1206 17798
rect 946 17412 970 17770
rect 1172 17412 1206 17770
rect 946 17386 1206 17412
rect 12370 17368 12400 18132
rect 12368 17290 12400 17368
rect 12502 17290 12540 18132
rect 23646 17930 24054 17976
rect 23646 17488 23674 17930
rect 24008 17488 24054 17930
rect 23646 17444 24054 17488
rect 12368 17240 12540 17290
rect 12368 17147 12534 17240
rect -313 16981 25321 17147
rect 11684 15874 13378 15926
rect 11736 13780 13362 13832
rect 11744 11696 13374 11748
rect 11720 9610 13416 9662
rect 11746 7524 13420 7576
rect 11726 5438 13352 5490
rect 11754 3354 13390 3406
rect 11662 1220 13430 1272
rect 19196 156 20478 188
rect 12470 108 12550 126
rect 4360 32 4916 94
rect 4360 -324 4412 32
rect 4854 -324 4916 32
rect 4360 -374 4916 -324
rect 12470 -472 12478 108
rect 12538 -472 12550 108
rect 19196 52 19222 156
rect 20440 52 20478 156
rect 19196 22 20478 52
rect 12470 -534 12550 -472
rect 12466 -568 12550 -534
rect 346 -652 25164 -568
rect 936 -788 1482 -688
rect 936 -1984 1006 -788
rect 1406 -1984 1482 -788
rect 8366 -744 8664 -698
rect 8366 -1102 8398 -744
rect 8632 -1102 8664 -744
rect 8366 -1446 8664 -1102
rect 16224 -750 16610 -706
rect 16224 -1082 16268 -750
rect 16572 -1082 16610 -750
rect 16224 -1464 16610 -1082
rect 23632 -752 24074 -694
rect 23632 -1826 23696 -752
rect 23998 -1826 24074 -752
rect 23632 -1902 24074 -1826
rect 936 -2064 1482 -1984
rect 6153 -2151 6219 -2008
<< via2 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 970 17412 1172 17770
rect 23674 17488 24008 17930
rect 4412 -324 4854 32
rect 19222 52 20440 156
rect 1006 -1984 1406 -788
rect 8398 -1102 8632 -744
rect 16268 -1082 16572 -750
rect 23696 -1826 23998 -752
<< metal3 >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
rect 23646 17970 24070 19418
rect 23502 17966 24070 17970
rect 15074 17930 24070 17966
rect 944 17770 10212 17800
rect 944 17412 970 17770
rect 1172 17412 10212 17770
rect 944 17280 10212 17412
rect 944 17276 1592 17280
rect 944 1099 1464 17276
rect 12066 15806 12180 17765
rect 12714 15813 12828 17841
rect 15074 17546 23674 17930
rect 23638 17488 23674 17546
rect 24008 17488 24070 17930
rect 23638 17444 24070 17488
rect 12910 15813 13417 15815
rect 11658 15805 12314 15806
rect 11658 15542 12400 15805
rect 12714 15573 13417 15813
rect 12714 15569 13244 15573
rect 11874 13734 12400 15542
rect 11674 13716 12400 13734
rect 11441 13470 12400 13716
rect 11874 11648 12400 13470
rect 11699 11402 12400 11648
rect 11874 9562 12400 11402
rect 11689 9316 12400 9562
rect 11874 7476 12400 9316
rect 11755 7230 12400 7476
rect 11874 5392 12400 7230
rect 11724 5146 12400 5392
rect 11874 3308 12400 5146
rect 11741 3062 12400 3308
rect 11874 1156 12400 3062
rect 944 1062 2019 1099
rect 944 1010 2033 1062
rect 11569 1026 12400 1156
rect 12718 13724 13244 15569
rect 12718 13478 13477 13724
rect 12718 11638 13244 13478
rect 12718 11392 13403 11638
rect 12718 9552 13244 11392
rect 12718 9306 13389 9552
rect 12718 7466 13244 9306
rect 12718 7220 13407 7466
rect 12718 5382 13244 7220
rect 12718 5136 13455 5382
rect 12718 1186 13244 5136
rect 944 1009 2019 1010
rect 944 -788 1464 1009
rect 11569 910 12402 1026
rect 12718 940 13523 1186
rect 23638 1120 24060 17444
rect 22984 1020 24060 1120
rect 12718 935 13244 940
rect 9784 698 10172 704
rect 9690 154 10172 698
rect 4360 32 4916 94
rect 4360 -324 4412 32
rect 4854 -324 4916 32
rect 4360 -374 4916 -324
rect 944 -1984 1006 -788
rect 1406 -1984 1464 -788
rect 8368 -744 8662 -694
rect 8368 -1102 8398 -744
rect 8632 -1102 8662 -744
rect 8368 -1152 8662 -1102
rect 9690 -1442 10166 154
rect 12218 -71 12288 910
rect 12728 -26 12812 935
rect 14904 696 15172 840
rect 14872 684 15172 696
rect 14366 154 15172 684
rect 14904 -1610 15172 154
rect 19196 156 20478 188
rect 19196 52 19222 156
rect 20440 52 20478 156
rect 19196 22 20478 52
rect 16228 -750 16616 -710
rect 16228 -1082 16268 -750
rect 16572 -1082 16616 -750
rect 16228 -1130 16616 -1082
rect 23638 -752 24060 1020
rect 23638 -1809 23696 -752
rect 944 -2052 1464 -1984
rect 20096 -1826 23696 -1809
rect 23998 -1826 24060 -752
rect 944 -2572 5348 -2052
rect 20096 -2231 24060 -1826
<< via3 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 4412 -324 4854 32
rect 8398 -1102 8632 -744
rect 19222 52 20440 156
rect 16268 -1082 16572 -750
<< metal4 >>
rect 649 22179 11573 22765
rect 649 12201 1235 22179
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
rect 9294 16326 15970 16902
rect 9306 14234 15754 14788
rect 667 128 1235 12201
rect 9346 12142 15794 12696
rect 9274 10042 15722 10596
rect 9200 7982 16026 8526
rect 9170 5872 15996 6416
rect 9170 3802 15996 4346
rect 9222 1670 16048 2214
rect 19196 156 20478 188
rect 4366 32 4904 100
rect 4366 -324 4412 32
rect 4854 -324 4904 32
rect 19196 52 19222 156
rect 20440 52 20478 156
rect 19196 22 20478 52
rect 4366 -2044 4904 -324
rect 8366 -744 8664 -698
rect 8366 -1102 8398 -744
rect 8632 -1102 8664 -744
rect 8366 -1446 8664 -1102
rect 16224 -750 16610 -706
rect 16224 -1082 16268 -750
rect 16572 -1082 16610 -750
rect 16224 -1464 16610 -1082
rect 20062 -1924 20474 22
rect 20630 -2014 20996 -2008
<< via4 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
<< metal5 >>
rect 13895 22499 25055 23089
rect 24465 18861 25055 22499
rect 18057 18772 25055 18861
rect 3340 18625 7634 18650
rect 0 18612 7634 18625
rect 0 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 25055 18772
rect 18057 18271 25055 18340
rect 0 18086 7634 18152
rect 0 18035 4377 18086
rect 0 14570 590 18035
rect 24465 16895 25055 18271
rect 9370 14854 16046 15430
rect 24465 14828 25083 16895
rect -8 14161 590 14570
rect -12 12853 590 14161
rect -12 12459 582 12853
rect 9294 12748 15742 13302
rect -12 11503 578 12459
rect -32 10235 578 11503
rect 9190 10658 15638 11212
rect -32 9379 558 10235
rect -32 798 572 9379
rect 9096 8568 15922 9112
rect 9054 6498 15880 7042
rect 9138 4408 15964 4952
rect 9138 2328 15964 2872
rect -32 194 2598 798
rect 24493 792 25083 14828
rect 9138 206 15964 750
rect 22598 232 25083 792
rect 22598 204 23864 232
use capacitor_8  capacitor_8_0
timestamp 1698679508
transform 1 0 1274 0 1 190
box 0 -430 10546 2050
use capacitor_8  capacitor_8_1
timestamp 1698679508
transform -1 0 23730 0 1 220
box 0 -430 10546 2050
use capacitors_1  capacitors_1_0
timestamp 1698684236
transform 1 0 1295 0 1 14846
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_1
timestamp 1698684236
transform -1 0 23807 0 1 14836
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_2
timestamp 1698684236
transform 1 0 1265 0 1 12742
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_3
timestamp 1698684236
transform 1 0 1269 0 1 10658
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_4
timestamp 1698684236
transform -1 0 23799 0 1 12752
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_5
timestamp 1698684236
transform -1 0 23775 0 1 10666
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_6
timestamp 1698684236
transform 1 0 1261 0 1 8572
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_7
timestamp 1698684236
transform 1 0 1251 0 1 6486
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_8
timestamp 1698684236
transform 1 0 1251 0 1 4400
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_9
timestamp 1698684236
transform 1 0 1263 0 1 2316
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_10
timestamp 1698684236
transform -1 0 23705 0 1 2296
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_11
timestamp 1698684236
transform -1 0 23727 0 1 4382
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_12
timestamp 1698684236
transform -1 0 23791 0 1 6466
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_13
timestamp 1698684236
transform -1 0 23831 0 1 8556
box -1291 -848 10655 2058
use clock  clock_0
timestamp 1698410772
transform 0 -1 12504 -1 0 25482
box -410 -1832 6030 1274
use nmos_dnw3  nmos_dnw3_0
timestamp 1698467949
transform 1 0 12184 0 1 16340
box -424 892 1176 2258
use pmos_cp1  pmos_cp1_0
timestamp 1698464655
transform 1 0 12196 0 -1 182
box -14 -278 858 754
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_0
timestamp 1698571947
transform -1 0 15980 0 1 -2156
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_1
timestamp 1698571947
transform 1 0 9038 0 1 -2176
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_2
timestamp 1698571947
transform 1 0 5164 0 1 -2412
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_3
timestamp 1698571947
transform -1 0 20174 0 1 -2456
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_4
timestamp 1698571947
transform -1 0 10140 0 1 18192
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_5
timestamp 1698571947
transform 1 0 15220 0 1 18184
box -1086 -940 1086 940
<< labels >>
rlabel metal3 12088 15446 12088 15446 1 input1
port 34 n
rlabel metal3 12964 15418 12964 15418 1 input2
port 35 n
rlabel metal4 964 12774 964 12774 1 vdd
port 1 n
rlabel metal5 24900 1146 24900 1146 1 gnd
port 64 n
rlabel metal2 12444 15904 12444 15904 1 in1
port 65 n
rlabel metal2 12576 11714 12576 11714 1 in3
port 66 n
rlabel metal2 12554 13796 12554 13796 1 in2
port 67 n
rlabel metal2 12598 9632 12598 9632 1 in4
port 68 n
rlabel metal2 12574 7544 12574 7544 1 in5
port 69 n
rlabel metal2 12526 5464 12526 5464 1 in6
port 70 n
rlabel metal2 12506 3382 12506 3382 1 in7
port 71 n
rlabel metal2 12554 1244 12554 1244 1 in8
port 73 n
<< end >>
