magic
tech sky130A
magscale 1 2
timestamp 1698683060
<< nwell >>
rect 44586 -1178 45022 -802
rect 50354 -1172 50790 -796
rect 67586 -1178 68022 -802
rect 73354 -1172 73790 -796
rect 91586 -1178 92022 -802
rect 97354 -1172 97790 -796
<< nmos >>
rect 44680 -1330 44710 -1246
rect 44898 -1330 44928 -1246
rect 50448 -1324 50478 -1240
rect 50666 -1324 50696 -1240
rect 67680 -1330 67710 -1246
rect 67898 -1330 67928 -1246
rect 73448 -1324 73478 -1240
rect 73666 -1324 73696 -1240
rect 91680 -1330 91710 -1246
rect 91898 -1330 91928 -1246
rect 97448 -1324 97478 -1240
rect 97666 -1324 97696 -1240
<< pmos >>
rect 44680 -1116 44710 -864
rect 44898 -1116 44928 -864
rect 50448 -1110 50478 -858
rect 50666 -1110 50696 -858
rect 67680 -1116 67710 -864
rect 67898 -1116 67928 -864
rect 73448 -1110 73478 -858
rect 73666 -1110 73696 -858
rect 91680 -1116 91710 -864
rect 91898 -1116 91928 -864
rect 97448 -1110 97478 -858
rect 97666 -1110 97696 -858
<< ndiff >>
rect 44622 -1258 44680 -1246
rect 44622 -1318 44634 -1258
rect 44668 -1318 44680 -1258
rect 44622 -1330 44680 -1318
rect 44710 -1258 44768 -1246
rect 44710 -1318 44722 -1258
rect 44756 -1318 44768 -1258
rect 44710 -1330 44768 -1318
rect 44840 -1258 44898 -1246
rect 44840 -1318 44852 -1258
rect 44886 -1318 44898 -1258
rect 44840 -1330 44898 -1318
rect 44928 -1258 44986 -1246
rect 44928 -1318 44940 -1258
rect 44974 -1318 44986 -1258
rect 44928 -1330 44986 -1318
rect 50390 -1252 50448 -1240
rect 50390 -1312 50402 -1252
rect 50436 -1312 50448 -1252
rect 50390 -1324 50448 -1312
rect 50478 -1252 50536 -1240
rect 50478 -1312 50490 -1252
rect 50524 -1312 50536 -1252
rect 50478 -1324 50536 -1312
rect 50608 -1252 50666 -1240
rect 50608 -1312 50620 -1252
rect 50654 -1312 50666 -1252
rect 50608 -1324 50666 -1312
rect 50696 -1252 50754 -1240
rect 50696 -1312 50708 -1252
rect 50742 -1312 50754 -1252
rect 50696 -1324 50754 -1312
rect 67622 -1258 67680 -1246
rect 67622 -1318 67634 -1258
rect 67668 -1318 67680 -1258
rect 67622 -1330 67680 -1318
rect 67710 -1258 67768 -1246
rect 67710 -1318 67722 -1258
rect 67756 -1318 67768 -1258
rect 67710 -1330 67768 -1318
rect 67840 -1258 67898 -1246
rect 67840 -1318 67852 -1258
rect 67886 -1318 67898 -1258
rect 67840 -1330 67898 -1318
rect 67928 -1258 67986 -1246
rect 67928 -1318 67940 -1258
rect 67974 -1318 67986 -1258
rect 67928 -1330 67986 -1318
rect 73390 -1252 73448 -1240
rect 73390 -1312 73402 -1252
rect 73436 -1312 73448 -1252
rect 73390 -1324 73448 -1312
rect 73478 -1252 73536 -1240
rect 73478 -1312 73490 -1252
rect 73524 -1312 73536 -1252
rect 73478 -1324 73536 -1312
rect 73608 -1252 73666 -1240
rect 73608 -1312 73620 -1252
rect 73654 -1312 73666 -1252
rect 73608 -1324 73666 -1312
rect 73696 -1252 73754 -1240
rect 73696 -1312 73708 -1252
rect 73742 -1312 73754 -1252
rect 73696 -1324 73754 -1312
rect 91622 -1258 91680 -1246
rect 91622 -1318 91634 -1258
rect 91668 -1318 91680 -1258
rect 91622 -1330 91680 -1318
rect 91710 -1258 91768 -1246
rect 91710 -1318 91722 -1258
rect 91756 -1318 91768 -1258
rect 91710 -1330 91768 -1318
rect 91840 -1258 91898 -1246
rect 91840 -1318 91852 -1258
rect 91886 -1318 91898 -1258
rect 91840 -1330 91898 -1318
rect 91928 -1258 91986 -1246
rect 91928 -1318 91940 -1258
rect 91974 -1318 91986 -1258
rect 91928 -1330 91986 -1318
rect 97390 -1252 97448 -1240
rect 97390 -1312 97402 -1252
rect 97436 -1312 97448 -1252
rect 97390 -1324 97448 -1312
rect 97478 -1252 97536 -1240
rect 97478 -1312 97490 -1252
rect 97524 -1312 97536 -1252
rect 97478 -1324 97536 -1312
rect 97608 -1252 97666 -1240
rect 97608 -1312 97620 -1252
rect 97654 -1312 97666 -1252
rect 97608 -1324 97666 -1312
rect 97696 -1252 97754 -1240
rect 97696 -1312 97708 -1252
rect 97742 -1312 97754 -1252
rect 97696 -1324 97754 -1312
<< pdiff >>
rect 44622 -876 44680 -864
rect 44622 -1104 44634 -876
rect 44668 -1104 44680 -876
rect 44622 -1116 44680 -1104
rect 44710 -876 44768 -864
rect 44710 -1104 44722 -876
rect 44756 -1104 44768 -876
rect 44710 -1116 44768 -1104
rect 44840 -876 44898 -864
rect 44840 -1104 44852 -876
rect 44886 -1104 44898 -876
rect 44840 -1116 44898 -1104
rect 44928 -876 44986 -864
rect 44928 -1104 44940 -876
rect 44974 -1104 44986 -876
rect 44928 -1116 44986 -1104
rect 50390 -870 50448 -858
rect 50390 -1098 50402 -870
rect 50436 -1098 50448 -870
rect 50390 -1110 50448 -1098
rect 50478 -870 50536 -858
rect 50478 -1098 50490 -870
rect 50524 -1098 50536 -870
rect 50478 -1110 50536 -1098
rect 50608 -870 50666 -858
rect 50608 -1098 50620 -870
rect 50654 -1098 50666 -870
rect 50608 -1110 50666 -1098
rect 50696 -870 50754 -858
rect 50696 -1098 50708 -870
rect 50742 -1098 50754 -870
rect 50696 -1110 50754 -1098
rect 67622 -876 67680 -864
rect 67622 -1104 67634 -876
rect 67668 -1104 67680 -876
rect 67622 -1116 67680 -1104
rect 67710 -876 67768 -864
rect 67710 -1104 67722 -876
rect 67756 -1104 67768 -876
rect 67710 -1116 67768 -1104
rect 67840 -876 67898 -864
rect 67840 -1104 67852 -876
rect 67886 -1104 67898 -876
rect 67840 -1116 67898 -1104
rect 67928 -876 67986 -864
rect 67928 -1104 67940 -876
rect 67974 -1104 67986 -876
rect 67928 -1116 67986 -1104
rect 73390 -870 73448 -858
rect 73390 -1098 73402 -870
rect 73436 -1098 73448 -870
rect 73390 -1110 73448 -1098
rect 73478 -870 73536 -858
rect 73478 -1098 73490 -870
rect 73524 -1098 73536 -870
rect 73478 -1110 73536 -1098
rect 73608 -870 73666 -858
rect 73608 -1098 73620 -870
rect 73654 -1098 73666 -870
rect 73608 -1110 73666 -1098
rect 73696 -870 73754 -858
rect 73696 -1098 73708 -870
rect 73742 -1098 73754 -870
rect 73696 -1110 73754 -1098
rect 91622 -876 91680 -864
rect 91622 -1104 91634 -876
rect 91668 -1104 91680 -876
rect 91622 -1116 91680 -1104
rect 91710 -876 91768 -864
rect 91710 -1104 91722 -876
rect 91756 -1104 91768 -876
rect 91710 -1116 91768 -1104
rect 91840 -876 91898 -864
rect 91840 -1104 91852 -876
rect 91886 -1104 91898 -876
rect 91840 -1116 91898 -1104
rect 91928 -876 91986 -864
rect 91928 -1104 91940 -876
rect 91974 -1104 91986 -876
rect 91928 -1116 91986 -1104
rect 97390 -870 97448 -858
rect 97390 -1098 97402 -870
rect 97436 -1098 97448 -870
rect 97390 -1110 97448 -1098
rect 97478 -870 97536 -858
rect 97478 -1098 97490 -870
rect 97524 -1098 97536 -870
rect 97478 -1110 97536 -1098
rect 97608 -870 97666 -858
rect 97608 -1098 97620 -870
rect 97654 -1098 97666 -870
rect 97608 -1110 97666 -1098
rect 97696 -870 97754 -858
rect 97696 -1098 97708 -870
rect 97742 -1098 97754 -870
rect 97696 -1110 97754 -1098
<< ndiffc >>
rect 44634 -1318 44668 -1258
rect 44722 -1318 44756 -1258
rect 44852 -1318 44886 -1258
rect 44940 -1318 44974 -1258
rect 50402 -1312 50436 -1252
rect 50490 -1312 50524 -1252
rect 50620 -1312 50654 -1252
rect 50708 -1312 50742 -1252
rect 67634 -1318 67668 -1258
rect 67722 -1318 67756 -1258
rect 67852 -1318 67886 -1258
rect 67940 -1318 67974 -1258
rect 73402 -1312 73436 -1252
rect 73490 -1312 73524 -1252
rect 73620 -1312 73654 -1252
rect 73708 -1312 73742 -1252
rect 91634 -1318 91668 -1258
rect 91722 -1318 91756 -1258
rect 91852 -1318 91886 -1258
rect 91940 -1318 91974 -1258
rect 97402 -1312 97436 -1252
rect 97490 -1312 97524 -1252
rect 97620 -1312 97654 -1252
rect 97708 -1312 97742 -1252
<< pdiffc >>
rect 44634 -1104 44668 -876
rect 44722 -1104 44756 -876
rect 44852 -1104 44886 -876
rect 44940 -1104 44974 -876
rect 50402 -1098 50436 -870
rect 50490 -1098 50524 -870
rect 50620 -1098 50654 -870
rect 50708 -1098 50742 -870
rect 67634 -1104 67668 -876
rect 67722 -1104 67756 -876
rect 67852 -1104 67886 -876
rect 67940 -1104 67974 -876
rect 73402 -1098 73436 -870
rect 73490 -1098 73524 -870
rect 73620 -1098 73654 -870
rect 73708 -1098 73742 -870
rect 91634 -1104 91668 -876
rect 91722 -1104 91756 -876
rect 91852 -1104 91886 -876
rect 91940 -1104 91974 -876
rect 97402 -1098 97436 -870
rect 97490 -1098 97524 -870
rect 97620 -1098 97654 -870
rect 97708 -1098 97742 -870
<< poly >>
rect 44680 -864 44710 -838
rect 44898 -864 44928 -838
rect 50448 -858 50478 -832
rect 50666 -858 50696 -832
rect 67680 -864 67710 -838
rect 67898 -864 67928 -838
rect 73448 -858 73478 -832
rect 73666 -858 73696 -832
rect 44362 -1172 44594 -1156
rect 44362 -1212 44380 -1172
rect 44574 -1174 44594 -1172
rect 44680 -1174 44710 -1116
rect 44898 -1154 44928 -1116
rect 44574 -1206 44710 -1174
rect 44574 -1212 44594 -1206
rect 44362 -1228 44594 -1212
rect 44680 -1246 44710 -1206
rect 44752 -1164 44928 -1154
rect 44752 -1200 44776 -1164
rect 44878 -1200 44928 -1164
rect 44752 -1210 44928 -1200
rect 44898 -1246 44928 -1210
rect 50130 -1166 50362 -1150
rect 50130 -1206 50148 -1166
rect 50342 -1168 50362 -1166
rect 50448 -1168 50478 -1110
rect 50666 -1148 50696 -1110
rect 91680 -864 91710 -838
rect 91898 -864 91928 -838
rect 97448 -858 97478 -832
rect 97666 -858 97696 -832
rect 50342 -1200 50478 -1168
rect 50342 -1206 50362 -1200
rect 50130 -1222 50362 -1206
rect 50448 -1240 50478 -1200
rect 50520 -1158 50696 -1148
rect 50520 -1194 50544 -1158
rect 50646 -1194 50696 -1158
rect 50520 -1204 50696 -1194
rect 50666 -1240 50696 -1204
rect 67362 -1172 67594 -1156
rect 67362 -1212 67380 -1172
rect 67574 -1174 67594 -1172
rect 67680 -1174 67710 -1116
rect 67898 -1154 67928 -1116
rect 67574 -1206 67710 -1174
rect 67574 -1212 67594 -1206
rect 67362 -1228 67594 -1212
rect 67680 -1246 67710 -1206
rect 67752 -1164 67928 -1154
rect 67752 -1200 67776 -1164
rect 67878 -1200 67928 -1164
rect 67752 -1210 67928 -1200
rect 67898 -1246 67928 -1210
rect 73130 -1166 73362 -1150
rect 73130 -1206 73148 -1166
rect 73342 -1168 73362 -1166
rect 73448 -1168 73478 -1110
rect 73666 -1148 73696 -1110
rect 73342 -1200 73478 -1168
rect 73342 -1206 73362 -1200
rect 73130 -1222 73362 -1206
rect 73448 -1240 73478 -1200
rect 73520 -1158 73696 -1148
rect 73520 -1194 73544 -1158
rect 73646 -1194 73696 -1158
rect 73520 -1204 73696 -1194
rect 73666 -1240 73696 -1204
rect 91362 -1172 91594 -1156
rect 91362 -1212 91380 -1172
rect 91574 -1174 91594 -1172
rect 91680 -1174 91710 -1116
rect 91898 -1154 91928 -1116
rect 91574 -1206 91710 -1174
rect 91574 -1212 91594 -1206
rect 91362 -1228 91594 -1212
rect 44680 -1356 44710 -1330
rect 44898 -1356 44928 -1330
rect 50448 -1350 50478 -1324
rect 50666 -1350 50696 -1324
rect 91680 -1246 91710 -1206
rect 91752 -1164 91928 -1154
rect 91752 -1200 91776 -1164
rect 91878 -1200 91928 -1164
rect 91752 -1210 91928 -1200
rect 91898 -1246 91928 -1210
rect 97130 -1166 97362 -1150
rect 97130 -1206 97148 -1166
rect 97342 -1168 97362 -1166
rect 97448 -1168 97478 -1110
rect 97666 -1148 97696 -1110
rect 97342 -1200 97478 -1168
rect 97342 -1206 97362 -1200
rect 97130 -1222 97362 -1206
rect 97448 -1240 97478 -1200
rect 97520 -1158 97696 -1148
rect 97520 -1194 97544 -1158
rect 97646 -1194 97696 -1158
rect 97520 -1204 97696 -1194
rect 97666 -1240 97696 -1204
rect 67680 -1356 67710 -1330
rect 67898 -1356 67928 -1330
rect 73448 -1350 73478 -1324
rect 73666 -1350 73696 -1324
rect 91680 -1356 91710 -1330
rect 91898 -1356 91928 -1330
rect 97448 -1350 97478 -1324
rect 97666 -1350 97696 -1324
<< polycont >>
rect 44380 -1212 44574 -1172
rect 44776 -1200 44878 -1164
rect 50148 -1206 50342 -1166
rect 50544 -1194 50646 -1158
rect 67380 -1212 67574 -1172
rect 67776 -1200 67878 -1164
rect 73148 -1206 73342 -1166
rect 73544 -1194 73646 -1158
rect 91380 -1212 91574 -1172
rect 91776 -1200 91878 -1164
rect 97148 -1206 97342 -1166
rect 97544 -1194 97646 -1158
<< locali >>
rect 44634 -876 44668 -860
rect 44634 -1120 44668 -1104
rect 44722 -876 44756 -860
rect 44722 -1120 44756 -1104
rect 44852 -876 44886 -860
rect 44852 -1120 44886 -1104
rect 44940 -876 44974 -860
rect 44940 -1120 44974 -1104
rect 50402 -870 50436 -854
rect 50402 -1114 50436 -1098
rect 50490 -870 50524 -854
rect 50490 -1114 50524 -1098
rect 50620 -870 50654 -854
rect 50620 -1114 50654 -1098
rect 50708 -870 50742 -854
rect 50708 -1114 50742 -1098
rect 67634 -876 67668 -860
rect 67634 -1120 67668 -1104
rect 67722 -876 67756 -860
rect 67722 -1120 67756 -1104
rect 67852 -876 67886 -860
rect 67852 -1120 67886 -1104
rect 67940 -876 67974 -860
rect 67940 -1120 67974 -1104
rect 73402 -870 73436 -854
rect 73402 -1114 73436 -1098
rect 73490 -870 73524 -854
rect 73490 -1114 73524 -1098
rect 73620 -870 73654 -854
rect 73620 -1114 73654 -1098
rect 73708 -870 73742 -854
rect 73708 -1114 73742 -1098
rect 91634 -876 91668 -860
rect 91634 -1120 91668 -1104
rect 91722 -876 91756 -860
rect 91722 -1120 91756 -1104
rect 91852 -876 91886 -860
rect 91852 -1120 91886 -1104
rect 91940 -876 91974 -860
rect 91940 -1120 91974 -1104
rect 97402 -870 97436 -854
rect 97402 -1114 97436 -1098
rect 97490 -870 97524 -854
rect 97490 -1114 97524 -1098
rect 97620 -870 97654 -854
rect 97620 -1114 97654 -1098
rect 97708 -870 97742 -854
rect 97708 -1114 97742 -1098
rect 44362 -1172 44594 -1156
rect 44362 -1212 44380 -1172
rect 44574 -1212 44594 -1172
rect 44752 -1164 44910 -1154
rect 44752 -1200 44776 -1164
rect 44878 -1200 44910 -1164
rect 44752 -1208 44910 -1200
rect 50130 -1166 50362 -1150
rect 50130 -1206 50148 -1166
rect 50342 -1206 50362 -1166
rect 50520 -1158 50678 -1148
rect 50520 -1194 50544 -1158
rect 50646 -1194 50678 -1158
rect 50520 -1202 50678 -1194
rect 44362 -1228 44594 -1212
rect 50130 -1222 50362 -1206
rect 67362 -1172 67594 -1156
rect 67362 -1212 67380 -1172
rect 67574 -1212 67594 -1172
rect 67752 -1164 67910 -1154
rect 67752 -1200 67776 -1164
rect 67878 -1200 67910 -1164
rect 67752 -1208 67910 -1200
rect 73130 -1166 73362 -1150
rect 73130 -1206 73148 -1166
rect 73342 -1206 73362 -1166
rect 73520 -1158 73678 -1148
rect 73520 -1194 73544 -1158
rect 73646 -1194 73678 -1158
rect 73520 -1202 73678 -1194
rect 67362 -1228 67594 -1212
rect 73130 -1222 73362 -1206
rect 91362 -1172 91594 -1156
rect 91362 -1212 91380 -1172
rect 91574 -1212 91594 -1172
rect 91752 -1164 91910 -1154
rect 91752 -1200 91776 -1164
rect 91878 -1200 91910 -1164
rect 91752 -1208 91910 -1200
rect 97130 -1166 97362 -1150
rect 97130 -1206 97148 -1166
rect 97342 -1206 97362 -1166
rect 97520 -1158 97678 -1148
rect 97520 -1194 97544 -1158
rect 97646 -1194 97678 -1158
rect 97520 -1202 97678 -1194
rect 91362 -1228 91594 -1212
rect 97130 -1222 97362 -1206
rect 44634 -1258 44668 -1242
rect 44634 -1334 44668 -1318
rect 44722 -1258 44756 -1242
rect 44722 -1334 44756 -1318
rect 44852 -1258 44886 -1242
rect 44852 -1334 44886 -1318
rect 44940 -1258 44974 -1242
rect 44940 -1334 44974 -1318
rect 50402 -1252 50436 -1236
rect 50402 -1328 50436 -1312
rect 50490 -1252 50524 -1236
rect 50490 -1328 50524 -1312
rect 50620 -1252 50654 -1236
rect 50620 -1328 50654 -1312
rect 50708 -1252 50742 -1236
rect 50708 -1328 50742 -1312
rect 67634 -1258 67668 -1242
rect 67634 -1334 67668 -1318
rect 67722 -1258 67756 -1242
rect 67722 -1334 67756 -1318
rect 67852 -1258 67886 -1242
rect 67852 -1334 67886 -1318
rect 67940 -1258 67974 -1242
rect 67940 -1334 67974 -1318
rect 73402 -1252 73436 -1236
rect 73402 -1328 73436 -1312
rect 73490 -1252 73524 -1236
rect 73490 -1328 73524 -1312
rect 73620 -1252 73654 -1236
rect 73620 -1328 73654 -1312
rect 73708 -1252 73742 -1236
rect 73708 -1328 73742 -1312
rect 91634 -1258 91668 -1242
rect 91634 -1334 91668 -1318
rect 91722 -1258 91756 -1242
rect 91722 -1334 91756 -1318
rect 91852 -1258 91886 -1242
rect 91852 -1334 91886 -1318
rect 91940 -1258 91974 -1242
rect 91940 -1334 91974 -1318
rect 97402 -1252 97436 -1236
rect 97402 -1328 97436 -1312
rect 97490 -1252 97524 -1236
rect 97490 -1328 97524 -1312
rect 97620 -1252 97654 -1236
rect 97620 -1328 97654 -1312
rect 97708 -1252 97742 -1236
rect 97708 -1328 97742 -1312
<< viali >>
rect 44634 -1104 44668 -876
rect 44722 -1104 44756 -876
rect 44852 -1104 44886 -876
rect 44940 -1104 44974 -876
rect 50402 -1098 50436 -870
rect 50490 -1098 50524 -870
rect 50620 -1098 50654 -870
rect 50708 -1098 50742 -870
rect 67634 -1104 67668 -876
rect 67722 -1104 67756 -876
rect 67852 -1104 67886 -876
rect 67940 -1104 67974 -876
rect 73402 -1098 73436 -870
rect 73490 -1098 73524 -870
rect 73620 -1098 73654 -870
rect 73708 -1098 73742 -870
rect 91634 -1104 91668 -876
rect 91722 -1104 91756 -876
rect 91852 -1104 91886 -876
rect 91940 -1104 91974 -876
rect 97402 -1098 97436 -870
rect 97490 -1098 97524 -870
rect 97620 -1098 97654 -870
rect 97708 -1098 97742 -870
rect 27274 -1214 27478 -1170
rect 44380 -1212 44574 -1172
rect 44776 -1200 44878 -1164
rect 50148 -1206 50342 -1166
rect 50544 -1194 50646 -1158
rect 51274 -1214 51478 -1170
rect 67380 -1212 67574 -1172
rect 67776 -1200 67878 -1164
rect 73148 -1206 73342 -1166
rect 73544 -1194 73646 -1158
rect 74274 -1214 74478 -1170
rect 91380 -1212 91574 -1172
rect 91776 -1200 91878 -1164
rect 97148 -1206 97342 -1166
rect 97544 -1194 97646 -1158
rect 98274 -1214 98478 -1170
rect 44634 -1318 44668 -1258
rect 44722 -1318 44756 -1258
rect 44852 -1318 44886 -1258
rect 44940 -1318 44974 -1258
rect 50402 -1312 50436 -1252
rect 50490 -1312 50524 -1252
rect 50620 -1312 50654 -1252
rect 50708 -1312 50742 -1252
rect 67634 -1318 67668 -1258
rect 67722 -1318 67756 -1258
rect 67852 -1318 67886 -1258
rect 67940 -1318 67974 -1258
rect 73402 -1312 73436 -1252
rect 73490 -1312 73524 -1252
rect 73620 -1312 73654 -1252
rect 73708 -1312 73742 -1252
rect 91634 -1318 91668 -1258
rect 91722 -1318 91756 -1258
rect 91852 -1318 91886 -1258
rect 91940 -1318 91974 -1258
rect 97402 -1312 97436 -1252
rect 97490 -1312 97524 -1252
rect 97620 -1312 97654 -1252
rect 97708 -1312 97742 -1252
<< metal1 >>
rect 44634 -816 44887 -782
rect 50402 -810 50655 -776
rect 44634 -864 44668 -816
rect 44852 -864 44886 -816
rect 50402 -858 50436 -810
rect 50620 -858 50654 -810
rect 67634 -816 67887 -782
rect 73402 -810 73655 -776
rect 44628 -876 44674 -864
rect 44628 -1104 44634 -876
rect 44668 -1104 44674 -876
rect 44628 -1116 44674 -1104
rect 44716 -876 44762 -864
rect 44716 -1104 44722 -876
rect 44756 -1104 44762 -876
rect 44716 -1116 44762 -1104
rect 44846 -876 44892 -864
rect 44846 -1104 44852 -876
rect 44886 -1104 44892 -876
rect 44846 -1116 44892 -1104
rect 44934 -876 44980 -864
rect 44934 -1104 44940 -876
rect 44974 -1104 44980 -876
rect 44934 -1116 44980 -1104
rect 50396 -870 50442 -858
rect 50396 -1098 50402 -870
rect 50436 -1098 50442 -870
rect 50396 -1110 50442 -1098
rect 50484 -870 50530 -858
rect 50484 -1098 50490 -870
rect 50524 -1098 50530 -870
rect 50484 -1110 50530 -1098
rect 50614 -870 50660 -858
rect 50614 -1098 50620 -870
rect 50654 -1098 50660 -870
rect 50614 -1110 50660 -1098
rect 50702 -870 50748 -858
rect 67634 -864 67668 -816
rect 67852 -864 67886 -816
rect 73402 -858 73436 -810
rect 73620 -858 73654 -810
rect 91634 -816 91887 -782
rect 97402 -810 97655 -776
rect 50702 -1098 50708 -870
rect 50742 -1098 50748 -870
rect 50702 -1110 50748 -1098
rect 67628 -876 67674 -864
rect 67628 -1104 67634 -876
rect 67668 -1104 67674 -876
rect 20940 -1176 26150 -1150
rect 44722 -1154 44756 -1116
rect 44940 -1150 44974 -1116
rect 50490 -1148 50524 -1110
rect 26742 -1170 27508 -1160
rect 26742 -1172 27274 -1170
rect 27478 -1172 27508 -1170
rect 20940 -1204 26338 -1176
rect 20940 -1218 26150 -1204
rect 26742 -1210 27268 -1172
rect 21010 -1222 26150 -1218
rect 27256 -1232 27268 -1210
rect 27490 -1232 27508 -1172
rect 44362 -1164 44594 -1156
rect 44362 -1222 44380 -1164
rect 44574 -1222 44594 -1164
rect 44362 -1228 44594 -1222
rect 44722 -1164 44910 -1154
rect 44722 -1200 44776 -1164
rect 44878 -1200 44910 -1164
rect 44722 -1210 44910 -1200
rect 44940 -1158 50362 -1150
rect 27256 -1242 27508 -1232
rect 44722 -1246 44756 -1210
rect 44940 -1216 50148 -1158
rect 50342 -1216 50362 -1158
rect 44940 -1218 50362 -1216
rect 44940 -1246 44974 -1218
rect 45010 -1222 50362 -1218
rect 50490 -1158 50678 -1148
rect 50490 -1194 50544 -1158
rect 50646 -1194 50678 -1158
rect 50490 -1204 50678 -1194
rect 50708 -1160 50742 -1110
rect 67628 -1116 67674 -1104
rect 67716 -876 67762 -864
rect 67716 -1104 67722 -876
rect 67756 -1104 67762 -876
rect 67716 -1116 67762 -1104
rect 67846 -876 67892 -864
rect 67846 -1104 67852 -876
rect 67886 -1104 67892 -876
rect 67846 -1116 67892 -1104
rect 67934 -876 67980 -864
rect 67934 -1104 67940 -876
rect 67974 -1104 67980 -876
rect 67934 -1116 67980 -1104
rect 73396 -870 73442 -858
rect 73396 -1098 73402 -870
rect 73436 -1098 73442 -870
rect 73396 -1110 73442 -1098
rect 73484 -870 73530 -858
rect 73484 -1098 73490 -870
rect 73524 -1098 73530 -870
rect 73484 -1110 73530 -1098
rect 73614 -870 73660 -858
rect 73614 -1098 73620 -870
rect 73654 -1098 73660 -870
rect 73614 -1110 73660 -1098
rect 73702 -870 73748 -858
rect 91634 -864 91668 -816
rect 91852 -864 91886 -816
rect 97402 -858 97436 -810
rect 97620 -858 97654 -810
rect 73702 -1098 73708 -870
rect 73742 -1098 73748 -870
rect 73702 -1110 73748 -1098
rect 91628 -876 91674 -864
rect 91628 -1104 91634 -876
rect 91668 -1104 91674 -876
rect 67722 -1154 67756 -1116
rect 67940 -1150 67974 -1116
rect 73490 -1148 73524 -1110
rect 50708 -1170 51508 -1160
rect 50708 -1172 51274 -1170
rect 51478 -1172 51508 -1170
rect 50490 -1240 50524 -1204
rect 50708 -1210 51268 -1172
rect 50708 -1240 50742 -1210
rect 51256 -1232 51268 -1210
rect 51490 -1232 51508 -1172
rect 67362 -1164 67594 -1156
rect 67362 -1222 67380 -1164
rect 67574 -1222 67594 -1164
rect 67362 -1228 67594 -1222
rect 67722 -1164 67910 -1154
rect 67722 -1200 67776 -1164
rect 67878 -1200 67910 -1164
rect 67722 -1210 67910 -1200
rect 67940 -1158 73362 -1150
rect 44628 -1258 44674 -1246
rect 44628 -1318 44634 -1258
rect 44668 -1318 44674 -1258
rect 44628 -1330 44674 -1318
rect 44716 -1258 44762 -1246
rect 44716 -1318 44722 -1258
rect 44756 -1318 44762 -1258
rect 44716 -1330 44762 -1318
rect 44846 -1258 44892 -1246
rect 44846 -1318 44852 -1258
rect 44886 -1318 44892 -1258
rect 44846 -1330 44892 -1318
rect 44934 -1258 44980 -1246
rect 44934 -1318 44940 -1258
rect 44974 -1318 44980 -1258
rect 44934 -1330 44980 -1318
rect 50396 -1252 50442 -1240
rect 50396 -1312 50402 -1252
rect 50436 -1312 50442 -1252
rect 50396 -1324 50442 -1312
rect 50484 -1252 50530 -1240
rect 50484 -1312 50490 -1252
rect 50524 -1312 50530 -1252
rect 50484 -1324 50530 -1312
rect 50614 -1252 50660 -1240
rect 50614 -1312 50620 -1252
rect 50654 -1312 50660 -1252
rect 50614 -1324 50660 -1312
rect 50702 -1252 50748 -1240
rect 51256 -1242 51508 -1232
rect 67722 -1246 67756 -1210
rect 67940 -1216 73148 -1158
rect 73342 -1216 73362 -1158
rect 67940 -1218 73362 -1216
rect 67940 -1246 67974 -1218
rect 68010 -1222 73362 -1218
rect 73490 -1158 73678 -1148
rect 73490 -1194 73544 -1158
rect 73646 -1194 73678 -1158
rect 73490 -1204 73678 -1194
rect 73708 -1160 73742 -1110
rect 91628 -1116 91674 -1104
rect 91716 -876 91762 -864
rect 91716 -1104 91722 -876
rect 91756 -1104 91762 -876
rect 91716 -1116 91762 -1104
rect 91846 -876 91892 -864
rect 91846 -1104 91852 -876
rect 91886 -1104 91892 -876
rect 91846 -1116 91892 -1104
rect 91934 -876 91980 -864
rect 91934 -1104 91940 -876
rect 91974 -1104 91980 -876
rect 91934 -1116 91980 -1104
rect 97396 -870 97442 -858
rect 97396 -1098 97402 -870
rect 97436 -1098 97442 -870
rect 97396 -1110 97442 -1098
rect 97484 -870 97530 -858
rect 97484 -1098 97490 -870
rect 97524 -1098 97530 -870
rect 97484 -1110 97530 -1098
rect 97614 -870 97660 -858
rect 97614 -1098 97620 -870
rect 97654 -1098 97660 -870
rect 97614 -1110 97660 -1098
rect 97702 -870 97748 -858
rect 97702 -1098 97708 -870
rect 97742 -1098 97748 -870
rect 97702 -1110 97748 -1098
rect 91722 -1154 91756 -1116
rect 91940 -1150 91974 -1116
rect 97490 -1148 97524 -1110
rect 73708 -1170 74508 -1160
rect 73708 -1172 74274 -1170
rect 74478 -1172 74508 -1170
rect 73490 -1240 73524 -1204
rect 73708 -1210 74268 -1172
rect 73708 -1240 73742 -1210
rect 74256 -1232 74268 -1210
rect 74490 -1232 74508 -1172
rect 91362 -1164 91594 -1156
rect 91362 -1222 91380 -1164
rect 91574 -1222 91594 -1164
rect 91362 -1228 91594 -1222
rect 91722 -1164 91910 -1154
rect 91722 -1200 91776 -1164
rect 91878 -1200 91910 -1164
rect 91722 -1210 91910 -1200
rect 91940 -1158 97362 -1150
rect 50702 -1312 50708 -1252
rect 50742 -1312 50748 -1252
rect 50702 -1324 50748 -1312
rect 67628 -1258 67674 -1246
rect 67628 -1318 67634 -1258
rect 67668 -1318 67674 -1258
rect 44634 -1358 44668 -1330
rect 44852 -1358 44886 -1330
rect 50402 -1352 50436 -1324
rect 50620 -1352 50654 -1324
rect 67628 -1330 67674 -1318
rect 67716 -1258 67762 -1246
rect 67716 -1318 67722 -1258
rect 67756 -1318 67762 -1258
rect 67716 -1330 67762 -1318
rect 67846 -1258 67892 -1246
rect 67846 -1318 67852 -1258
rect 67886 -1318 67892 -1258
rect 67846 -1330 67892 -1318
rect 67934 -1258 67980 -1246
rect 67934 -1318 67940 -1258
rect 67974 -1318 67980 -1258
rect 67934 -1330 67980 -1318
rect 73396 -1252 73442 -1240
rect 73396 -1312 73402 -1252
rect 73436 -1312 73442 -1252
rect 73396 -1324 73442 -1312
rect 73484 -1252 73530 -1240
rect 73484 -1312 73490 -1252
rect 73524 -1312 73530 -1252
rect 73484 -1324 73530 -1312
rect 73614 -1252 73660 -1240
rect 73614 -1312 73620 -1252
rect 73654 -1312 73660 -1252
rect 73614 -1324 73660 -1312
rect 73702 -1252 73748 -1240
rect 74256 -1242 74508 -1232
rect 91722 -1246 91756 -1210
rect 91940 -1216 97148 -1158
rect 97342 -1216 97362 -1158
rect 91940 -1218 97362 -1216
rect 91940 -1246 91974 -1218
rect 92010 -1222 97362 -1218
rect 97490 -1158 97678 -1148
rect 97490 -1194 97544 -1158
rect 97646 -1194 97678 -1158
rect 97490 -1204 97678 -1194
rect 97708 -1160 97742 -1110
rect 97708 -1170 98508 -1160
rect 97708 -1172 98274 -1170
rect 98478 -1172 98508 -1170
rect 97490 -1240 97524 -1204
rect 97708 -1210 98268 -1172
rect 97708 -1240 97742 -1210
rect 98256 -1232 98268 -1210
rect 98490 -1232 98508 -1172
rect 73702 -1312 73708 -1252
rect 73742 -1312 73748 -1252
rect 73702 -1324 73748 -1312
rect 91628 -1258 91674 -1246
rect 91628 -1318 91634 -1258
rect 91668 -1318 91674 -1258
rect 67634 -1358 67668 -1330
rect 67852 -1358 67886 -1330
rect 73402 -1352 73436 -1324
rect 73620 -1352 73654 -1324
rect 91628 -1330 91674 -1318
rect 91716 -1258 91762 -1246
rect 91716 -1318 91722 -1258
rect 91756 -1318 91762 -1258
rect 91716 -1330 91762 -1318
rect 91846 -1258 91892 -1246
rect 91846 -1318 91852 -1258
rect 91886 -1318 91892 -1258
rect 91846 -1330 91892 -1318
rect 91934 -1258 91980 -1246
rect 91934 -1318 91940 -1258
rect 91974 -1318 91980 -1258
rect 91934 -1330 91980 -1318
rect 97396 -1252 97442 -1240
rect 97396 -1312 97402 -1252
rect 97436 -1312 97442 -1252
rect 97396 -1324 97442 -1312
rect 97484 -1252 97530 -1240
rect 97484 -1312 97490 -1252
rect 97524 -1312 97530 -1252
rect 97484 -1324 97530 -1312
rect 97614 -1252 97660 -1240
rect 97614 -1312 97620 -1252
rect 97654 -1312 97660 -1252
rect 97614 -1324 97660 -1312
rect 97702 -1252 97748 -1240
rect 98256 -1242 98508 -1232
rect 97702 -1312 97708 -1252
rect 97742 -1312 97748 -1252
rect 97702 -1324 97748 -1312
rect 91634 -1358 91668 -1330
rect 91852 -1358 91886 -1330
rect 97402 -1352 97436 -1324
rect 97620 -1352 97654 -1324
<< via1 >>
rect 27268 -1214 27274 -1172
rect 27274 -1214 27478 -1172
rect 27478 -1214 27490 -1172
rect 27268 -1232 27490 -1214
rect 44380 -1172 44574 -1164
rect 44380 -1212 44574 -1172
rect 44380 -1222 44574 -1212
rect 50148 -1166 50342 -1158
rect 50148 -1206 50342 -1166
rect 50148 -1216 50342 -1206
rect 51268 -1214 51274 -1172
rect 51274 -1214 51478 -1172
rect 51478 -1214 51490 -1172
rect 51268 -1232 51490 -1214
rect 67380 -1172 67574 -1164
rect 67380 -1212 67574 -1172
rect 67380 -1222 67574 -1212
rect 73148 -1166 73342 -1158
rect 73148 -1206 73342 -1166
rect 73148 -1216 73342 -1206
rect 74268 -1214 74274 -1172
rect 74274 -1214 74478 -1172
rect 74478 -1214 74490 -1172
rect 74268 -1232 74490 -1214
rect 91380 -1172 91574 -1164
rect 91380 -1212 91574 -1172
rect 91380 -1222 91574 -1212
rect 97148 -1166 97342 -1158
rect 97148 -1206 97342 -1166
rect 97148 -1216 97342 -1206
rect 98268 -1214 98274 -1172
rect 98274 -1214 98478 -1172
rect 98478 -1214 98490 -1172
rect 98268 -1232 98490 -1214
<< metal2 >>
rect 44480 25420 46872 25660
rect 46632 24910 46872 25420
rect 91012 25410 94204 25650
rect 93964 24900 94204 25410
rect -108 23650 1682 23730
rect 25044 23722 25284 23734
rect 21716 23660 25284 23722
rect 45020 23670 48556 23726
rect 68452 23672 71968 23732
rect 25044 23594 25284 23660
rect 91694 23658 95834 23720
rect -16 21560 1774 21640
rect 21738 21584 25270 21646
rect 45036 21578 48572 21634
rect 68438 21574 71954 21634
rect 91682 21576 95822 21638
rect 21710 19618 21884 19626
rect 21710 19566 21916 19618
rect 36 19468 1826 19548
rect 21710 19510 25350 19566
rect 21728 19482 25350 19510
rect 45028 19492 48564 19548
rect 68426 19482 71942 19542
rect 91690 19482 95830 19544
rect 21636 17470 21828 17502
rect 102 17378 1892 17458
rect 21636 17442 25294 17470
rect 21636 17386 25328 17442
rect 45018 17406 48554 17462
rect 68360 17400 71876 17460
rect 91690 17386 95830 17448
rect 25056 17328 25328 17386
rect 50 15278 1840 15358
rect 21662 15314 25284 15398
rect 45020 15304 48556 15360
rect 68350 15302 71866 15362
rect 91686 15288 95826 15350
rect 128 13200 1918 13280
rect 21636 13224 25186 13270
rect 45102 13208 48610 13278
rect 68358 13218 71874 13278
rect 91774 13212 95914 13274
rect 132 11106 1922 11186
rect 21742 11118 25124 11190
rect 45096 11114 48604 11184
rect 68358 11120 71874 11180
rect 91760 11118 95900 11180
rect 126 9020 1916 9100
rect 21678 9032 25060 9104
rect 45096 9026 48604 9096
rect 68358 9026 71854 9106
rect 91764 9020 95904 9082
rect 23392 7344 23572 7974
rect 69950 7346 70190 7952
rect 11784 7104 23578 7344
rect 67368 7106 70190 7346
rect 20374 -1160 20574 -1150
rect 44374 -1156 44574 -1150
rect 44362 -1160 44594 -1156
rect 20374 -1228 20574 -1218
rect 27268 -1172 27490 -1162
rect 44362 -1218 44374 -1160
rect 44362 -1222 44380 -1218
rect 44574 -1222 44594 -1160
rect 50130 -1158 50362 -1150
rect 67374 -1156 67574 -1150
rect 50130 -1216 50148 -1158
rect 50342 -1216 50362 -1158
rect 67362 -1160 67594 -1156
rect 50130 -1222 50362 -1216
rect 51268 -1172 51490 -1162
rect 44362 -1228 44594 -1222
rect 27268 -1242 27490 -1232
rect 67362 -1218 67374 -1160
rect 67362 -1222 67380 -1218
rect 67574 -1222 67594 -1160
rect 73130 -1158 73362 -1150
rect 91374 -1156 91574 -1150
rect 73130 -1216 73148 -1158
rect 73342 -1216 73362 -1158
rect 91362 -1160 91594 -1156
rect 73130 -1222 73362 -1216
rect 74268 -1172 74490 -1162
rect 67362 -1228 67594 -1222
rect 51268 -1242 51490 -1232
rect 91362 -1218 91374 -1160
rect 91362 -1222 91380 -1218
rect 91574 -1222 91594 -1160
rect 97130 -1158 97362 -1150
rect 97130 -1216 97148 -1158
rect 97342 -1216 97362 -1158
rect 97130 -1222 97362 -1216
rect 98268 -1172 98490 -1162
rect 91362 -1228 91594 -1222
rect 74268 -1242 74490 -1232
rect 98268 -1242 98490 -1232
<< via2 >>
rect 20374 -1218 20574 -1160
rect 27268 -1232 27490 -1172
rect 44374 -1164 44574 -1160
rect 44374 -1218 44380 -1164
rect 44380 -1218 44574 -1164
rect 51268 -1232 51490 -1172
rect 67374 -1164 67574 -1160
rect 67374 -1218 67380 -1164
rect 67380 -1218 67574 -1164
rect 74268 -1232 74490 -1172
rect 91374 -1164 91574 -1160
rect 91374 -1218 91380 -1164
rect 91380 -1218 91574 -1164
rect 98268 -1232 98490 -1172
<< metal3 >>
rect 11892 -1760 11964 294
rect 20208 -1155 20570 -1148
rect 20208 -1160 20584 -1155
rect 20208 -1216 20374 -1160
rect 20212 -1740 20280 -1216
rect 20364 -1218 20374 -1216
rect 20574 -1218 20584 -1160
rect 20364 -1223 20584 -1218
rect 27258 -1170 27500 -1167
rect 27258 -1172 28032 -1170
rect 27258 -1232 27268 -1172
rect 27490 -1232 28032 -1172
rect 27258 -1237 28032 -1232
rect 27270 -1242 28032 -1237
rect 17014 -1760 17084 -1756
rect 20212 -1760 20274 -1740
rect -417 -2314 20274 -1760
rect 11892 -2320 11964 -2314
rect 17014 -2315 17084 -2314
rect 20212 -2316 20274 -2314
rect 27954 -1760 28026 -1242
rect 34918 -1760 34990 -766
rect 44208 -1155 44570 -1148
rect 44208 -1160 44584 -1155
rect 44208 -1216 44374 -1160
rect 44212 -1358 44280 -1216
rect 44364 -1218 44374 -1216
rect 44574 -1218 44584 -1160
rect 44364 -1223 44584 -1218
rect 51258 -1170 51500 -1167
rect 51258 -1172 52032 -1170
rect 51258 -1232 51268 -1172
rect 51490 -1232 52032 -1172
rect 51258 -1237 52032 -1232
rect 51270 -1242 52032 -1237
rect 44212 -1760 44278 -1358
rect 51954 -1760 52026 -1242
rect 58636 -1760 58708 296
rect 67208 -1155 67570 -1148
rect 91208 -1155 91570 -1148
rect 67208 -1160 67584 -1155
rect 67208 -1216 67374 -1160
rect 67212 -1358 67280 -1216
rect 67364 -1218 67374 -1216
rect 67574 -1218 67584 -1160
rect 91208 -1160 91584 -1155
rect 67364 -1223 67584 -1218
rect 74258 -1170 74500 -1167
rect 74258 -1172 75032 -1170
rect 74258 -1232 74268 -1172
rect 74490 -1232 75032 -1172
rect 91208 -1216 91374 -1160
rect 74258 -1237 75032 -1232
rect 74270 -1242 75032 -1237
rect 67212 -1760 67278 -1358
rect 74954 -1760 75026 -1242
rect 91212 -1358 91280 -1216
rect 91364 -1218 91374 -1216
rect 91574 -1218 91584 -1160
rect 91364 -1223 91584 -1218
rect 98258 -1170 98500 -1167
rect 98258 -1172 99032 -1170
rect 98258 -1232 98268 -1172
rect 98490 -1232 99032 -1172
rect 98258 -1237 99032 -1232
rect 98270 -1242 99032 -1237
rect 91212 -1760 91278 -1358
rect 98954 -1760 99026 -1242
rect 27954 -2314 44278 -1760
rect 51952 -2314 67278 -1760
rect 74952 -2314 91282 -1760
rect 98948 -2314 117458 -1760
rect 27954 -2322 28026 -2314
rect 51954 -2316 52026 -2314
rect 58636 -2318 58708 -2314
rect 67212 -2315 67278 -2314
rect 91212 -2315 91278 -2314
<< metal4 >>
rect 878 -2703 1536 3251
rect 41173 -2703 41831 2795
rect 52613 2513 54547 3171
rect 53303 -2703 53961 2513
rect 87553 -2703 88211 2769
rect 100311 -2703 100969 3147
rect 878 -3361 100969 -2703
<< metal5 >>
rect 284 -3683 942 8622
rect 29877 -3683 30535 2977
rect 63777 -3683 64435 3163
rect 78167 -3683 78825 2967
rect 116571 -3683 117161 4223
rect 284 -4341 117170 -3683
rect 284 -4350 942 -4341
rect 116571 -4359 117161 -4341
use buffer_digital  buffer_digital_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698389822
transform 1 0 20636 0 1 -1358
box -274 0 412 576
use buffer_digital  buffer_digital_1
timestamp 1698389822
transform 1 0 26404 0 1 -1352
box -274 0 412 576
use charge_pump  charge_pump_0 ~/Desktop/charge_pumps2/layout_files2
timestamp 1698675553
transform 1 0 -480 0 1 7870
box 498 -7862 23756 19014
use charge_pump  charge_pump_1
timestamp 1698675553
transform 1 0 46226 0 1 7872
box 498 -7862 23756 19014
use charge_pump  charge_pump_2
timestamp 1698675553
transform 1 0 93528 0 1 7864
box 498 -7862 23756 19014
use charge_pump_reverse  charge_pump_reverse_0 ~/Desktop/charge_pumps2/layout_files2
timestamp 1698672105
transform 1 0 22894 0 -1 24894
box 498 -3206 23756 25968
use charge_pump_reverse  charge_pump_reverse_1
timestamp 1698672105
transform 1 0 69556 0 -1 24884
box 498 -3206 23756 25968
<< end >>
