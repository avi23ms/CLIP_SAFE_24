magic
tech sky130A
magscale 1 2
timestamp 1698873245
<< error_p >>
rect -29 551 29 557
rect -29 517 -17 551
rect -29 511 29 517
rect -29 311 29 317
rect -29 277 -17 311
rect -29 271 29 277
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -169 29 -163
rect -29 -203 -17 -169
rect -29 -209 29 -203
rect -29 -409 29 -403
rect -29 -443 -17 -409
rect -29 -449 29 -443
rect -29 -649 29 -643
rect -29 -683 -17 -649
rect -29 -689 29 -683
<< nmos >>
rect -15 589 15 673
rect -15 349 15 433
rect -15 109 15 193
rect -15 -131 15 -47
rect -15 -371 15 -287
rect -15 -611 15 -527
<< ndiff >>
rect -73 661 -15 673
rect -73 601 -61 661
rect -27 601 -15 661
rect -73 589 -15 601
rect 15 661 73 673
rect 15 601 27 661
rect 61 601 73 661
rect 15 589 73 601
rect -73 421 -15 433
rect -73 361 -61 421
rect -27 361 -15 421
rect -73 349 -15 361
rect 15 421 73 433
rect 15 361 27 421
rect 61 361 73 421
rect 15 349 73 361
rect -73 181 -15 193
rect -73 121 -61 181
rect -27 121 -15 181
rect -73 109 -15 121
rect 15 181 73 193
rect 15 121 27 181
rect 61 121 73 181
rect 15 109 73 121
rect -73 -59 -15 -47
rect -73 -119 -61 -59
rect -27 -119 -15 -59
rect -73 -131 -15 -119
rect 15 -59 73 -47
rect 15 -119 27 -59
rect 61 -119 73 -59
rect 15 -131 73 -119
rect -73 -299 -15 -287
rect -73 -359 -61 -299
rect -27 -359 -15 -299
rect -73 -371 -15 -359
rect 15 -299 73 -287
rect 15 -359 27 -299
rect 61 -359 73 -299
rect 15 -371 73 -359
rect -73 -539 -15 -527
rect -73 -599 -61 -539
rect -27 -599 -15 -539
rect -73 -611 -15 -599
rect 15 -539 73 -527
rect 15 -599 27 -539
rect 61 -599 73 -539
rect 15 -611 73 -599
<< ndiffc >>
rect -61 601 -27 661
rect 27 601 61 661
rect -61 361 -27 421
rect 27 361 61 421
rect -61 121 -27 181
rect 27 121 61 181
rect -61 -119 -27 -59
rect 27 -119 61 -59
rect -61 -359 -27 -299
rect 27 -359 61 -299
rect -61 -599 -27 -539
rect 27 -599 61 -539
<< poly >>
rect -15 673 15 699
rect -15 567 15 589
rect -33 551 33 567
rect -33 517 -17 551
rect 17 517 33 551
rect -33 501 33 517
rect -15 433 15 459
rect -15 327 15 349
rect -33 311 33 327
rect -33 277 -17 311
rect 17 277 33 311
rect -33 261 33 277
rect -15 193 15 219
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -15 -47 15 -21
rect -15 -153 15 -131
rect -33 -169 33 -153
rect -33 -203 -17 -169
rect 17 -203 33 -169
rect -33 -219 33 -203
rect -15 -287 15 -261
rect -15 -393 15 -371
rect -33 -409 33 -393
rect -33 -443 -17 -409
rect 17 -443 33 -409
rect -33 -459 33 -443
rect -15 -527 15 -501
rect -15 -633 15 -611
rect -33 -649 33 -633
rect -33 -683 -17 -649
rect 17 -683 33 -649
rect -33 -699 33 -683
<< polycont >>
rect -17 517 17 551
rect -17 277 17 311
rect -17 37 17 71
rect -17 -203 17 -169
rect -17 -443 17 -409
rect -17 -683 17 -649
<< locali >>
rect -61 661 -27 677
rect -61 585 -27 601
rect 27 661 61 677
rect 27 585 61 601
rect -33 517 -17 551
rect 17 517 33 551
rect -61 421 -27 437
rect -61 345 -27 361
rect 27 421 61 437
rect 27 345 61 361
rect -33 277 -17 311
rect 17 277 33 311
rect -61 181 -27 197
rect -61 105 -27 121
rect 27 181 61 197
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -61 -59 -27 -43
rect -61 -135 -27 -119
rect 27 -59 61 -43
rect 27 -135 61 -119
rect -33 -203 -17 -169
rect 17 -203 33 -169
rect -61 -299 -27 -283
rect -61 -375 -27 -359
rect 27 -299 61 -283
rect 27 -375 61 -359
rect -33 -443 -17 -409
rect 17 -443 33 -409
rect -61 -539 -27 -523
rect -61 -615 -27 -599
rect 27 -539 61 -523
rect 27 -615 61 -599
rect -33 -683 -17 -649
rect 17 -683 33 -649
<< viali >>
rect -61 601 -27 661
rect 27 601 61 661
rect -17 517 17 551
rect -61 361 -27 421
rect 27 361 61 421
rect -17 277 17 311
rect -61 121 -27 181
rect 27 121 61 181
rect -17 37 17 71
rect -61 -119 -27 -59
rect 27 -119 61 -59
rect -17 -203 17 -169
rect -61 -359 -27 -299
rect 27 -359 61 -299
rect -17 -443 17 -409
rect -61 -599 -27 -539
rect 27 -599 61 -539
rect -17 -683 17 -649
<< metal1 >>
rect -67 661 -21 673
rect -67 601 -61 661
rect -27 601 -21 661
rect -67 589 -21 601
rect 21 661 67 673
rect 21 601 27 661
rect 61 601 67 661
rect 21 589 67 601
rect -29 551 29 557
rect -29 517 -17 551
rect 17 517 29 551
rect -29 511 29 517
rect -67 421 -21 433
rect -67 361 -61 421
rect -27 361 -21 421
rect -67 349 -21 361
rect 21 421 67 433
rect 21 361 27 421
rect 61 361 67 421
rect 21 349 67 361
rect -29 311 29 317
rect -29 277 -17 311
rect 17 277 29 311
rect -29 271 29 277
rect -67 181 -21 193
rect -67 121 -61 181
rect -27 121 -21 181
rect -67 109 -21 121
rect 21 181 67 193
rect 21 121 27 181
rect 61 121 67 181
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -67 -59 -21 -47
rect -67 -119 -61 -59
rect -27 -119 -21 -59
rect -67 -131 -21 -119
rect 21 -59 67 -47
rect 21 -119 27 -59
rect 61 -119 67 -59
rect 21 -131 67 -119
rect -29 -169 29 -163
rect -29 -203 -17 -169
rect 17 -203 29 -169
rect -29 -209 29 -203
rect -67 -299 -21 -287
rect -67 -359 -61 -299
rect -27 -359 -21 -299
rect -67 -371 -21 -359
rect 21 -299 67 -287
rect 21 -359 27 -299
rect 61 -359 67 -299
rect 21 -371 67 -359
rect -29 -409 29 -403
rect -29 -443 -17 -409
rect 17 -443 29 -409
rect -29 -449 29 -443
rect -67 -539 -21 -527
rect -67 -599 -61 -539
rect -27 -599 -21 -539
rect -67 -611 -21 -599
rect 21 -539 67 -527
rect 21 -599 27 -539
rect 61 -599 67 -539
rect 21 -611 67 -599
rect -29 -649 29 -643
rect -29 -683 -17 -649
rect 17 -683 29 -649
rect -29 -689 29 -683
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 6 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
