magic
tech sky130A
magscale 1 2
timestamp 1697915631
<< pwell >>
rect -641 -810 641 810
<< nmos >>
rect -445 -600 -345 600
rect -287 -600 -187 600
rect -129 -600 -29 600
rect 29 -600 129 600
rect 187 -600 287 600
rect 345 -600 445 600
<< ndiff >>
rect -503 588 -445 600
rect -503 -588 -491 588
rect -457 -588 -445 588
rect -503 -600 -445 -588
rect -345 588 -287 600
rect -345 -588 -333 588
rect -299 -588 -287 588
rect -345 -600 -287 -588
rect -187 588 -129 600
rect -187 -588 -175 588
rect -141 -588 -129 588
rect -187 -600 -129 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 129 588 187 600
rect 129 -588 141 588
rect 175 -588 187 588
rect 129 -600 187 -588
rect 287 588 345 600
rect 287 -588 299 588
rect 333 -588 345 588
rect 287 -600 345 -588
rect 445 588 503 600
rect 445 -588 457 588
rect 491 -588 503 588
rect 445 -600 503 -588
<< ndiffc >>
rect -491 -588 -457 588
rect -333 -588 -299 588
rect -175 -588 -141 588
rect -17 -588 17 588
rect 141 -588 175 588
rect 299 -588 333 588
rect 457 -588 491 588
<< psubdiff >>
rect -605 740 -509 774
rect 509 740 605 774
rect -605 678 -571 740
rect 571 678 605 740
rect -605 -740 -571 -678
rect 571 -740 605 -678
rect -605 -774 -509 -740
rect 509 -774 605 -740
<< psubdiffcont >>
rect -509 740 509 774
rect -605 -678 -571 678
rect 571 -678 605 678
rect -509 -774 509 -740
<< poly >>
rect -445 672 -345 688
rect -445 638 -429 672
rect -361 638 -345 672
rect -445 600 -345 638
rect -287 672 -187 688
rect -287 638 -271 672
rect -203 638 -187 672
rect -287 600 -187 638
rect -129 672 -29 688
rect -129 638 -113 672
rect -45 638 -29 672
rect -129 600 -29 638
rect 29 672 129 688
rect 29 638 45 672
rect 113 638 129 672
rect 29 600 129 638
rect 187 672 287 688
rect 187 638 203 672
rect 271 638 287 672
rect 187 600 287 638
rect 345 672 445 688
rect 345 638 361 672
rect 429 638 445 672
rect 345 600 445 638
rect -445 -638 -345 -600
rect -445 -672 -429 -638
rect -361 -672 -345 -638
rect -445 -688 -345 -672
rect -287 -638 -187 -600
rect -287 -672 -271 -638
rect -203 -672 -187 -638
rect -287 -688 -187 -672
rect -129 -638 -29 -600
rect -129 -672 -113 -638
rect -45 -672 -29 -638
rect -129 -688 -29 -672
rect 29 -638 129 -600
rect 29 -672 45 -638
rect 113 -672 129 -638
rect 29 -688 129 -672
rect 187 -638 287 -600
rect 187 -672 203 -638
rect 271 -672 287 -638
rect 187 -688 287 -672
rect 345 -638 445 -600
rect 345 -672 361 -638
rect 429 -672 445 -638
rect 345 -688 445 -672
<< polycont >>
rect -429 638 -361 672
rect -271 638 -203 672
rect -113 638 -45 672
rect 45 638 113 672
rect 203 638 271 672
rect 361 638 429 672
rect -429 -672 -361 -638
rect -271 -672 -203 -638
rect -113 -672 -45 -638
rect 45 -672 113 -638
rect 203 -672 271 -638
rect 361 -672 429 -638
<< locali >>
rect -605 740 -509 774
rect 509 740 605 774
rect -605 678 -571 740
rect 571 678 605 740
rect -445 638 -429 672
rect -361 638 -345 672
rect -287 638 -271 672
rect -203 638 -187 672
rect -129 638 -113 672
rect -45 638 -29 672
rect 29 638 45 672
rect 113 638 129 672
rect 187 638 203 672
rect 271 638 287 672
rect 345 638 361 672
rect 429 638 445 672
rect -491 588 -457 604
rect -491 -604 -457 -588
rect -333 588 -299 604
rect -333 -604 -299 -588
rect -175 588 -141 604
rect -175 -604 -141 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 141 588 175 604
rect 141 -604 175 -588
rect 299 588 333 604
rect 299 -604 333 -588
rect 457 588 491 604
rect 457 -604 491 -588
rect -445 -672 -429 -638
rect -361 -672 -345 -638
rect -287 -672 -271 -638
rect -203 -672 -187 -638
rect -129 -672 -113 -638
rect -45 -672 -29 -638
rect 29 -672 45 -638
rect 113 -672 129 -638
rect 187 -672 203 -638
rect 271 -672 287 -638
rect 345 -672 361 -638
rect 429 -672 445 -638
rect -605 -740 -571 -678
rect 571 -740 605 -678
rect -605 -774 -509 -740
rect 509 -774 605 -740
<< viali >>
rect -429 638 -361 672
rect -271 638 -203 672
rect -113 638 -45 672
rect 45 638 113 672
rect 203 638 271 672
rect 361 638 429 672
rect -491 -588 -457 588
rect -333 -588 -299 588
rect -175 -588 -141 588
rect -17 -588 17 588
rect 141 -588 175 588
rect 299 -588 333 588
rect 457 -588 491 588
rect -429 -672 -361 -638
rect -271 -672 -203 -638
rect -113 -672 -45 -638
rect 45 -672 113 -638
rect 203 -672 271 -638
rect 361 -672 429 -638
<< metal1 >>
rect -441 672 -349 678
rect -441 638 -429 672
rect -361 638 -349 672
rect -441 632 -349 638
rect -283 672 -191 678
rect -283 638 -271 672
rect -203 638 -191 672
rect -283 632 -191 638
rect -125 672 -33 678
rect -125 638 -113 672
rect -45 638 -33 672
rect -125 632 -33 638
rect 33 672 125 678
rect 33 638 45 672
rect 113 638 125 672
rect 33 632 125 638
rect 191 672 283 678
rect 191 638 203 672
rect 271 638 283 672
rect 191 632 283 638
rect 349 672 441 678
rect 349 638 361 672
rect 429 638 441 672
rect 349 632 441 638
rect -497 588 -451 600
rect -497 -588 -491 588
rect -457 -588 -451 588
rect -497 -600 -451 -588
rect -339 588 -293 600
rect -339 -588 -333 588
rect -299 -588 -293 588
rect -339 -600 -293 -588
rect -181 588 -135 600
rect -181 -588 -175 588
rect -141 -588 -135 588
rect -181 -600 -135 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 135 588 181 600
rect 135 -588 141 588
rect 175 -588 181 588
rect 135 -600 181 -588
rect 293 588 339 600
rect 293 -588 299 588
rect 333 -588 339 588
rect 293 -600 339 -588
rect 451 588 497 600
rect 451 -588 457 588
rect 491 -588 497 588
rect 451 -600 497 -588
rect -441 -638 -349 -632
rect -441 -672 -429 -638
rect -361 -672 -349 -638
rect -441 -678 -349 -672
rect -283 -638 -191 -632
rect -283 -672 -271 -638
rect -203 -672 -191 -638
rect -283 -678 -191 -672
rect -125 -638 -33 -632
rect -125 -672 -113 -638
rect -45 -672 -33 -638
rect -125 -678 -33 -672
rect 33 -638 125 -632
rect 33 -672 45 -638
rect 113 -672 125 -638
rect 33 -678 125 -672
rect 191 -638 283 -632
rect 191 -672 203 -638
rect 271 -672 283 -638
rect 191 -678 283 -672
rect 349 -638 441 -632
rect 349 -672 361 -638
rect 429 -672 441 -638
rect 349 -678 441 -672
<< properties >>
string FIXED_BBOX -588 -757 588 757
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6 l 0.5 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
