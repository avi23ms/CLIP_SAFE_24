magic
tech sky130A
magscale 1 2
timestamp 1698179620
<< metal1 >>
rect 150 1513 312 1583
rect 3226 1550 3236 1614
rect 3334 1550 3344 1614
rect 1788 970 1804 1002
rect 1878 982 1976 986
rect 1878 914 1914 982
rect 1986 914 1996 982
rect 1878 902 1976 914
rect 477 656 582 659
rect 470 604 480 656
rect 564 604 582 656
rect 3474 626 3540 662
rect 477 577 582 604
rect 3558 442 3912 490
rect 270 409 312 442
rect 2078 256 3731 266
rect 1064 230 3731 256
rect 1064 214 2132 230
rect 3654 172 3731 230
rect 3680 35 3731 172
rect 770 -129 813 -59
rect 2874 -66 2884 -42
rect 2498 -114 2884 -66
rect 2970 -114 2980 -42
rect 1764 -234 1826 -198
rect 1730 -348 1740 -286
rect 1712 -372 1740 -348
rect 1792 -372 1802 -286
rect 1712 -390 1776 -372
rect 1482 -780 1540 -752
rect 1780 -776 1838 -748
rect 3680 -966 3728 35
rect 3438 -1014 3728 -966
rect 3864 -1066 3912 442
rect 2491 -1126 2804 -1077
rect 3668 -1114 3912 -1066
<< via1 >>
rect 3236 1550 3334 1614
rect 1914 914 1986 982
rect 480 604 564 656
rect 2884 -114 2970 -42
rect 1740 -372 1792 -286
<< metal2 >>
rect 3236 1614 3334 1624
rect 3334 1556 3660 1611
rect 3236 1540 3334 1550
rect 1914 982 1986 992
rect 1986 924 2636 972
rect 1914 904 1986 914
rect 480 656 564 666
rect 480 594 564 604
rect 492 -1128 532 594
rect 880 14 920 872
rect 880 -26 1796 14
rect 1756 -276 1796 -26
rect 1740 -286 1796 -276
rect 1792 -372 1796 -286
rect 1740 -382 1792 -372
rect 2588 -430 2636 924
rect 2884 -42 2970 -32
rect 3605 -54 3660 1556
rect 2970 -106 3660 -54
rect 3605 -107 3660 -106
rect 2884 -124 2970 -114
rect 1808 -478 2636 -430
use cmfb  cmfb_0
timestamp 1698179620
transform 1 0 -54 0 1 -439
box 203 439 3639 2056
use integrator_new1  integrator_new1_0
timestamp 1698177474
transform 1 0 -1633 0 1 -3755
box 1247 441 5619 3693
<< labels >>
rlabel metal2 3641 577 3641 577 1 Vdd
port 1 n
rlabel metal1 3895 -938 3895 -938 1 gnd
port 2 n
rlabel metal1 1524 -768 1524 -768 1 vin1
port 3 n
rlabel metal1 1788 -767 1788 -767 1 vin2
port 4 n
rlabel metal1 1268 233 1268 233 1 Vbias
port 5 n
rlabel metal1 3513 647 3513 647 1 Vcmref
port 6 n
rlabel metal2 997 -14 997 -14 1 vo2
port 7 n
rlabel metal2 510 -659 510 -659 1 vo1
port 8 n
<< end >>
