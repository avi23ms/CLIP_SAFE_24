magic
tech sky130A
magscale 1 2
timestamp 1699103691
<< dnwell >>
rect -254 2098 880 2232
rect -324 2078 880 2098
rect -324 2048 1074 2078
rect -400 2034 1074 2048
rect -418 1130 1074 2034
rect -324 1086 1074 1130
rect -254 1070 1074 1086
rect -254 906 880 1070
<< nwell >>
rect 544 2256 1176 2258
rect -424 2040 1176 2256
rect -424 1130 -252 2040
rect 952 1130 1176 2040
rect -424 896 1176 1130
rect -194 894 1176 896
rect 512 892 1176 894
<< nmos >>
rect 94 1858 124 1942
rect 422 1858 452 1942
rect 4 1200 204 1800
rect 330 1200 530 1800
<< ndiff >>
rect 32 1928 94 1942
rect 32 1872 46 1928
rect 80 1872 94 1928
rect 32 1858 94 1872
rect 124 1920 184 1942
rect 124 1882 140 1920
rect 174 1882 184 1920
rect 124 1858 184 1882
rect 362 1920 422 1942
rect 362 1882 372 1920
rect 406 1882 422 1920
rect 362 1858 422 1882
rect 452 1928 514 1942
rect 452 1872 466 1928
rect 500 1872 514 1928
rect 452 1858 514 1872
rect -106 1770 4 1800
rect -106 1230 -76 1770
rect -26 1230 4 1770
rect -106 1200 4 1230
rect 204 1778 330 1800
rect 204 1230 234 1778
rect 296 1230 330 1778
rect 204 1200 330 1230
rect 530 1770 640 1800
rect 530 1230 560 1770
rect 610 1230 640 1770
rect 530 1200 640 1230
<< ndiffc >>
rect 46 1872 80 1928
rect 140 1882 174 1920
rect 372 1882 406 1920
rect 466 1872 500 1928
rect -76 1230 -26 1770
rect 234 1230 296 1778
rect 560 1230 610 1770
<< psubdiff >>
rect 828 1460 912 1496
rect 828 1286 850 1460
rect 894 1286 912 1460
rect 828 1250 912 1286
<< nsubdiff >>
rect 1018 1460 1102 1496
rect 1018 1286 1038 1460
rect 1082 1286 1102 1460
rect 1018 1250 1102 1286
<< psubdiffcont >>
rect 850 1286 894 1460
<< nsubdiffcont >>
rect 1038 1286 1082 1460
<< poly >>
rect 302 2138 452 2150
rect 302 2104 324 2138
rect 430 2104 452 2138
rect 302 2090 452 2104
rect 94 2054 248 2066
rect 94 2020 118 2054
rect 224 2020 248 2054
rect 94 2006 248 2020
rect 94 1942 124 2006
rect 422 1942 452 2090
rect 94 1826 124 1858
rect 422 1826 452 1858
rect 4 1800 204 1826
rect 330 1800 530 1826
rect 4 1172 204 1200
rect 330 1174 530 1200
<< polycont >>
rect 324 2104 430 2138
rect 118 2020 224 2054
<< locali >>
rect 302 2138 452 2150
rect 302 2104 324 2138
rect 430 2104 452 2138
rect 302 2090 452 2104
rect 94 2054 248 2066
rect 94 2020 118 2054
rect 224 2020 248 2054
rect 94 2006 248 2020
rect 34 1928 90 1944
rect 132 1936 182 1942
rect 34 1872 46 1928
rect 80 1872 90 1928
rect 34 1854 90 1872
rect 130 1924 184 1936
rect 130 1878 140 1924
rect 130 1864 184 1878
rect 366 1920 416 1946
rect 366 1882 372 1920
rect 406 1882 416 1920
rect 132 1856 182 1864
rect 366 1854 416 1882
rect 456 1928 512 1944
rect 456 1872 466 1928
rect 500 1872 512 1928
rect 456 1854 512 1872
rect -98 1770 2 1796
rect -98 1734 -76 1770
rect -26 1768 2 1770
rect -96 1230 -76 1734
rect -24 1734 2 1768
rect 206 1778 328 1818
rect 542 1790 640 1800
rect -24 1234 -6 1734
rect -26 1230 -6 1234
rect -96 1210 -6 1230
rect 206 1230 234 1778
rect 296 1230 328 1778
rect 206 1188 328 1230
rect 540 1770 640 1790
rect 540 1230 560 1770
rect 610 1766 640 1770
rect 612 1758 640 1766
rect 612 1234 630 1758
rect 828 1460 1102 1496
rect 828 1286 850 1460
rect 894 1286 1038 1460
rect 1082 1286 1102 1460
rect 828 1250 1102 1286
rect 610 1230 630 1234
rect 540 1210 630 1230
<< viali >>
rect 324 2104 430 2138
rect 118 2020 224 2054
rect 46 1872 80 1928
rect 140 1920 184 1924
rect 140 1882 174 1920
rect 174 1882 184 1920
rect 140 1878 184 1882
rect 372 1882 406 1920
rect 466 1872 500 1928
rect -76 1234 -26 1768
rect -26 1234 -24 1768
rect 234 1230 296 1778
rect 560 1234 610 1766
rect 610 1234 612 1766
<< metal1 >>
rect -78 2138 452 2150
rect -78 2104 324 2138
rect 430 2104 452 2138
rect -78 2094 452 2104
rect -78 1944 -22 2094
rect 304 2090 452 2094
rect 94 2062 248 2066
rect 94 2010 118 2062
rect 224 2010 248 2062
rect 94 2006 248 2010
rect 34 1944 90 1946
rect -152 1928 92 1944
rect 132 1936 182 1942
rect 366 1936 416 1946
rect -152 1872 46 1928
rect 80 1872 92 1928
rect -152 1856 92 1872
rect 130 1924 416 1936
rect 130 1878 140 1924
rect 184 1920 416 1924
rect 184 1882 372 1920
rect 406 1882 416 1920
rect 184 1878 416 1882
rect 130 1864 416 1878
rect 132 1856 326 1864
rect 34 1854 90 1856
rect 204 1818 326 1856
rect 366 1854 416 1864
rect 454 1938 698 1944
rect 454 1928 564 1938
rect 454 1872 466 1928
rect 500 1872 564 1928
rect 454 1860 564 1872
rect 636 1860 698 1938
rect 454 1856 698 1860
rect 456 1854 512 1856
rect -108 1772 4 1794
rect 204 1788 328 1818
rect -108 1230 -98 1772
rect -6 1230 4 1772
rect -108 1202 4 1230
rect 206 1778 328 1788
rect 206 1230 234 1778
rect 296 1230 328 1778
rect -96 1194 -6 1202
rect 206 1188 328 1230
rect 530 1772 640 1794
rect 530 1230 544 1772
rect 626 1269 640 1772
rect 626 1230 641 1269
rect 530 1202 641 1230
rect 551 1194 641 1202
<< via1 >>
rect 118 2054 224 2062
rect 118 2020 224 2054
rect 118 2010 224 2020
rect 564 1860 636 1938
rect -98 1768 -6 1772
rect -98 1234 -76 1768
rect -76 1234 -24 1768
rect -24 1234 -6 1768
rect -98 1230 -6 1234
rect 544 1766 626 1772
rect 544 1234 560 1766
rect 560 1234 612 1766
rect 612 1234 626 1766
rect 544 1230 626 1234
<< metal2 >>
rect 94 2062 644 2066
rect 94 2010 118 2062
rect 224 2010 644 2062
rect 94 2006 644 2010
rect 556 1938 644 2006
rect 556 1860 564 1938
rect 636 1860 644 1938
rect 556 1856 644 1860
rect -108 1772 4 1794
rect -108 1230 -98 1772
rect -6 1230 4 1772
rect -108 1202 4 1230
rect 530 1772 640 1794
rect 530 1230 544 1772
rect 626 1230 640 1772
rect 530 1202 640 1230
<< via2 >>
rect -98 1230 -6 1772
rect 544 1230 626 1772
<< metal3 >>
rect -108 1772 4 1794
rect -108 1230 -98 1772
rect -6 1230 4 1772
rect 530 1772 640 1794
rect 530 1268 544 1772
rect -108 1216 4 1230
rect 528 1230 544 1268
rect 626 1230 640 1772
rect 528 1204 640 1230
<< labels >>
rlabel metal1 254 1888 254 1888 1 vin
port 1 n
rlabel metal2 -52 1210 -52 1210 1 out1
port 2 n
rlabel metal3 590 1210 590 1210 1 out2
port 3 n
rlabel metal1 -66 1896 -66 1896 1 clk
port 4 n
rlabel metal1 680 1916 680 1916 1 clkb
port 5 n
rlabel nwell -372 1752 -372 1752 1 vs
port 6 n
<< end >>
