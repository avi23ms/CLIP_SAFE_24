magic
tech sky130A
magscale 1 2
timestamp 1698652801
<< nwell >>
rect -401 104 401 142
rect -497 -142 497 104
<< pmos >>
rect -399 -42 -369 42
rect -303 -42 -273 42
rect -207 -42 -177 42
rect -111 -42 -81 42
rect -15 -42 15 42
rect 81 -42 111 42
rect 177 -42 207 42
rect 273 -42 303 42
rect 369 -42 399 42
<< pdiff >>
rect -461 30 -399 42
rect -461 -30 -449 30
rect -415 -30 -399 30
rect -461 -42 -399 -30
rect -369 30 -303 42
rect -369 -30 -353 30
rect -319 -30 -303 30
rect -369 -42 -303 -30
rect -273 30 -207 42
rect -273 -30 -257 30
rect -223 -30 -207 30
rect -273 -42 -207 -30
rect -177 30 -111 42
rect -177 -30 -161 30
rect -127 -30 -111 30
rect -177 -42 -111 -30
rect -81 30 -15 42
rect -81 -30 -65 30
rect -31 -30 -15 30
rect -81 -42 -15 -30
rect 15 30 81 42
rect 15 -30 31 30
rect 65 -30 81 30
rect 15 -42 81 -30
rect 111 30 177 42
rect 111 -30 127 30
rect 161 -30 177 30
rect 111 -42 177 -30
rect 207 30 273 42
rect 207 -30 223 30
rect 257 -30 273 30
rect 207 -42 273 -30
rect 303 30 369 42
rect 303 -30 319 30
rect 353 -30 369 30
rect 303 -42 369 -30
rect 399 30 461 42
rect 399 -30 415 30
rect 449 -30 461 30
rect 399 -42 461 -30
<< pdiffc >>
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
<< poly >>
rect -321 123 -255 139
rect -321 89 -305 123
rect -271 89 -255 123
rect -321 73 -255 89
rect -129 123 -63 139
rect -129 89 -113 123
rect -79 89 -63 123
rect -129 73 -63 89
rect 63 123 129 139
rect 63 89 79 123
rect 113 89 129 123
rect 63 73 129 89
rect 255 123 321 139
rect 255 89 271 123
rect 305 89 321 123
rect 255 73 321 89
rect -399 42 -369 68
rect -303 42 -273 73
rect -207 42 -177 68
rect -111 42 -81 73
rect -15 42 15 68
rect 81 42 111 73
rect 177 42 207 68
rect 273 42 303 73
rect 369 42 399 68
rect -399 -73 -369 -42
rect -303 -68 -273 -42
rect -207 -73 -177 -42
rect -111 -68 -81 -42
rect -15 -73 15 -42
rect 81 -68 111 -42
rect 177 -73 207 -42
rect 273 -68 303 -42
rect 369 -73 399 -42
rect -417 -89 -351 -73
rect -417 -123 -401 -89
rect -367 -123 -351 -89
rect -417 -139 -351 -123
rect -225 -89 -159 -73
rect -225 -123 -209 -89
rect -175 -123 -159 -89
rect -225 -139 -159 -123
rect -33 -89 33 -73
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect -33 -139 33 -123
rect 159 -89 225 -73
rect 159 -123 175 -89
rect 209 -123 225 -89
rect 159 -139 225 -123
rect 351 -89 417 -73
rect 351 -123 367 -89
rect 401 -123 417 -89
rect 351 -139 417 -123
<< polycont >>
rect -305 89 -271 123
rect -113 89 -79 123
rect 79 89 113 123
rect 271 89 305 123
rect -401 -123 -367 -89
rect -209 -123 -175 -89
rect -17 -123 17 -89
rect 175 -123 209 -89
rect 367 -123 401 -89
<< locali >>
rect -321 89 -305 123
rect -271 89 -255 123
rect -129 89 -113 123
rect -79 89 -63 123
rect 63 89 79 123
rect 113 89 129 123
rect 255 89 271 123
rect 305 89 321 123
rect -449 30 -415 46
rect -449 -46 -415 -30
rect -353 30 -319 46
rect -353 -46 -319 -30
rect -257 30 -223 46
rect -257 -46 -223 -30
rect -161 30 -127 46
rect -161 -46 -127 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 127 30 161 46
rect 127 -46 161 -30
rect 223 30 257 46
rect 223 -46 257 -30
rect 319 30 353 46
rect 319 -46 353 -30
rect 415 30 449 46
rect 415 -46 449 -30
rect -417 -123 -401 -89
rect -367 -123 -351 -89
rect -225 -123 -209 -89
rect -175 -123 -159 -89
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect 159 -123 175 -89
rect 209 -123 225 -89
rect 351 -123 367 -89
rect 401 -123 417 -89
<< viali >>
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
<< metal1 >>
rect -455 30 -409 42
rect -455 -30 -449 30
rect -415 -30 -409 30
rect -455 -42 -409 -30
rect -359 30 -313 42
rect -359 -30 -353 30
rect -319 -30 -313 30
rect -359 -42 -313 -30
rect -263 30 -217 42
rect -263 -30 -257 30
rect -223 -30 -217 30
rect -263 -42 -217 -30
rect -167 30 -121 42
rect -167 -30 -161 30
rect -127 -30 -121 30
rect -167 -42 -121 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 121 30 167 42
rect 121 -30 127 30
rect 161 -30 167 30
rect 121 -42 167 -30
rect 217 30 263 42
rect 217 -30 223 30
rect 257 -30 263 30
rect 217 -42 263 -30
rect 313 30 359 42
rect 313 -30 319 30
rect 353 -30 359 30
rect 313 -42 359 -30
rect 409 30 455 42
rect 409 -30 415 30
rect 449 -30 455 30
rect 409 -42 455 -30
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 9 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
