magic
tech sky130A
magscale 1 2
timestamp 1698611618
<< error_p >>
rect -365 114 -307 120
rect -173 114 -115 120
rect 19 114 77 120
rect 211 114 269 120
rect 403 114 461 120
rect -365 80 -353 114
rect -173 80 -161 114
rect 19 80 31 114
rect 211 80 223 114
rect 403 80 415 114
rect -365 74 -307 80
rect -173 74 -115 80
rect 19 74 77 80
rect 211 74 269 80
rect 403 74 461 80
rect -461 -80 -403 -74
rect -269 -80 -211 -74
rect -77 -80 -19 -74
rect 115 -80 173 -74
rect 307 -80 365 -74
rect -461 -114 -449 -80
rect -269 -114 -257 -80
rect -77 -114 -65 -80
rect 115 -114 127 -80
rect 307 -114 319 -80
rect -461 -120 -403 -114
rect -269 -120 -211 -114
rect -77 -120 -19 -114
rect 115 -120 173 -114
rect 307 -120 365 -114
<< nmos >>
rect -447 -42 -417 42
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
rect 417 -42 447 42
<< ndiff >>
rect -509 30 -447 42
rect -509 -30 -497 30
rect -463 -30 -447 30
rect -509 -42 -447 -30
rect -417 30 -351 42
rect -417 -30 -401 30
rect -367 -30 -351 30
rect -417 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 417 42
rect 351 -30 367 30
rect 401 -30 417 30
rect 351 -42 417 -30
rect 447 30 509 42
rect 447 -30 463 30
rect 497 -30 509 30
rect 447 -42 509 -30
<< ndiffc >>
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
<< poly >>
rect -369 114 -303 130
rect -369 80 -353 114
rect -319 80 -303 114
rect -447 42 -417 68
rect -369 64 -303 80
rect -177 114 -111 130
rect -177 80 -161 114
rect -127 80 -111 114
rect -351 42 -321 64
rect -255 42 -225 68
rect -177 64 -111 80
rect 15 114 81 130
rect 15 80 31 114
rect 65 80 81 114
rect -159 42 -129 64
rect -63 42 -33 68
rect 15 64 81 80
rect 207 114 273 130
rect 207 80 223 114
rect 257 80 273 114
rect 33 42 63 64
rect 129 42 159 68
rect 207 64 273 80
rect 399 114 465 130
rect 399 80 415 114
rect 449 80 465 114
rect 225 42 255 64
rect 321 42 351 68
rect 399 64 465 80
rect 417 42 447 64
rect -447 -64 -417 -42
rect -465 -80 -399 -64
rect -351 -68 -321 -42
rect -255 -64 -225 -42
rect -465 -114 -449 -80
rect -415 -114 -399 -80
rect -465 -130 -399 -114
rect -273 -80 -207 -64
rect -159 -68 -129 -42
rect -63 -64 -33 -42
rect -273 -114 -257 -80
rect -223 -114 -207 -80
rect -273 -130 -207 -114
rect -81 -80 -15 -64
rect 33 -68 63 -42
rect 129 -64 159 -42
rect -81 -114 -65 -80
rect -31 -114 -15 -80
rect -81 -130 -15 -114
rect 111 -80 177 -64
rect 225 -68 255 -42
rect 321 -64 351 -42
rect 111 -114 127 -80
rect 161 -114 177 -80
rect 111 -130 177 -114
rect 303 -80 369 -64
rect 417 -68 447 -42
rect 303 -114 319 -80
rect 353 -114 369 -80
rect 303 -130 369 -114
<< polycont >>
rect -353 80 -319 114
rect -161 80 -127 114
rect 31 80 65 114
rect 223 80 257 114
rect 415 80 449 114
rect -449 -114 -415 -80
rect -257 -114 -223 -80
rect -65 -114 -31 -80
rect 127 -114 161 -80
rect 319 -114 353 -80
<< locali >>
rect -369 80 -353 114
rect -319 80 -303 114
rect -177 80 -161 114
rect -127 80 -111 114
rect 15 80 31 114
rect 65 80 81 114
rect 207 80 223 114
rect 257 80 273 114
rect 399 80 415 114
rect 449 80 465 114
rect -497 30 -463 46
rect -497 -46 -463 -30
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect 463 30 497 46
rect 463 -46 497 -30
rect -465 -114 -449 -80
rect -415 -114 -399 -80
rect -273 -114 -257 -80
rect -223 -114 -207 -80
rect -81 -114 -65 -80
rect -31 -114 -15 -80
rect 111 -114 127 -80
rect 161 -114 177 -80
rect 303 -114 319 -80
rect 353 -114 369 -80
<< viali >>
rect -353 80 -319 114
rect -161 80 -127 114
rect 31 80 65 114
rect 223 80 257 114
rect 415 80 449 114
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect -449 -114 -415 -80
rect -257 -114 -223 -80
rect -65 -114 -31 -80
rect 127 -114 161 -80
rect 319 -114 353 -80
<< metal1 >>
rect -365 114 -307 120
rect -365 80 -353 114
rect -319 80 -307 114
rect -365 74 -307 80
rect -173 114 -115 120
rect -173 80 -161 114
rect -127 80 -115 114
rect -173 74 -115 80
rect 19 114 77 120
rect 19 80 31 114
rect 65 80 77 114
rect 19 74 77 80
rect 211 114 269 120
rect 211 80 223 114
rect 257 80 269 114
rect 211 74 269 80
rect 403 114 461 120
rect 403 80 415 114
rect 449 80 461 114
rect 403 74 461 80
rect -503 30 -457 42
rect -503 -30 -497 30
rect -463 -30 -457 30
rect -503 -42 -457 -30
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect 457 30 503 42
rect 457 -30 463 30
rect 497 -30 503 30
rect 457 -42 503 -30
rect -461 -80 -403 -74
rect -461 -114 -449 -80
rect -415 -114 -403 -80
rect -461 -120 -403 -114
rect -269 -80 -211 -74
rect -269 -114 -257 -80
rect -223 -114 -211 -80
rect -269 -120 -211 -114
rect -77 -80 -19 -74
rect -77 -114 -65 -80
rect -31 -114 -19 -80
rect -77 -120 -19 -114
rect 115 -80 173 -74
rect 115 -114 127 -80
rect 161 -114 173 -80
rect 115 -120 173 -114
rect 307 -80 365 -74
rect 307 -114 319 -80
rect 353 -114 365 -80
rect 307 -120 365 -114
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
