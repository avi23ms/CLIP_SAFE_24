magic
tech sky130A
magscale 1 2
timestamp 1699130246
<< nwell >>
rect 228 1148 684 1466
rect 228 1094 704 1148
rect 866 1094 1238 1466
rect 228 1012 1238 1094
rect 1380 -364 3438 -124
rect 7118 -356 8214 -142
<< nsubdiff >>
rect 3296 -234 3402 -210
rect 3296 -298 3320 -234
rect 3378 -298 3402 -234
rect 3296 -316 3402 -298
rect 8064 -234 8174 -208
rect 8064 -290 8094 -234
rect 8146 -290 8174 -234
rect 8064 -318 8174 -290
<< nsubdiffcont >>
rect 3320 -298 3378 -234
rect 8094 -290 8146 -234
<< locali >>
rect 3296 -234 3402 -210
rect 3296 -298 3320 -234
rect 3378 -298 3402 -234
rect 3296 -316 3402 -298
rect 8070 -234 8176 -204
rect 8070 -290 8094 -234
rect 8146 -290 8176 -234
rect 8070 -318 8176 -290
<< viali >>
rect 3320 -298 3378 -234
rect 8094 -290 8146 -234
<< metal1 >>
rect 738 1478 862 1814
rect 742 528 858 548
rect 768 486 836 528
rect 3296 -234 3402 -210
rect 3296 -298 3320 -234
rect 3378 -298 3402 -234
rect 3296 -316 3402 -298
rect 7114 -234 8194 -202
rect 7114 -290 8094 -234
rect 8146 -290 8194 -234
rect 7114 -306 8194 -290
use capacito7  capacitor_7_0
timestamp 1699130246
transform 1 0 739 0 1 0
box -739 -430 9807 2050
<< end >>
