* SPICE3 file created from reconfigurable_CP_lvs1.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_1_MH6KF8 c1_n1046_n900# m3_n1086_n940# VSUBS
X0 c1_n1046_n900# m3_n1086_n940# sky130_fd_pr__cap_mim_m3_1 l=9 w=9
C0 m3_n1086_n940# c1_n1046_n900# 7.77654f
C1 m3_n1086_n940# VSUBS 3.30833f
.ends

.subckt sky130_fd_pr__pfet_01v8_FXZ64Q a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_DQBD8A a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt buffer_digital i in VDD GND a_116_148#
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 VDD VDD a_116_148# i GND sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 VDD VDD in a_116_148# GND sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 a_116_148# i GND GND sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 in a_116_148# GND GND sky130_fd_pr__nfet_01v8_DQBD8A
.ends

.subckt sky130_fd_pr__nfet_01v8_D4CMYK a_15_n130# a_63_n42# a_n177_n130# a_255_n42#
+ a_n129_n42# a_111_64# a_n321_n42# a_159_n42# a_n81_64# a_n273_64# a_351_n42# a_207_n130#
+ a_303_64# a_n33_n42# a_n369_n130# a_n225_n42# a_n413_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_n130# a_n413_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_4ZKXAA a_63_n42# a_n417_n42# a_303_n139# w_n545_n142#
+ a_255_n42# a_n465_n139# a_n129_n42# a_111_n139# a_447_n42# a_n273_n139# a_n177_73#
+ a_n321_n42# a_207_73# a_n509_n42# a_159_n42# a_15_73# a_n81_n139# a_351_n42# a_n33_n42#
+ a_n369_73# a_n225_n42# a_399_73# VSUBS
X0 a_n33_n42# a_n81_n139# a_n129_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_351_n42# a_303_n139# a_255_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n139# a_63_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_73# a_159_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_447_n42# a_399_73# a_351_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_73# a_n417_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n225_n42# a_n273_n139# a_n321_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n139# a_n509_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X8 a_n129_n42# a_n177_73# a_n225_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_63_n42# a_15_73# a_n33_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC45 a_63_n42# a_15_64# a_n417_n42# a_111_n130#
+ a_n273_n130# a_255_n42# a_n129_n42# a_n369_64# a_399_64# a_447_n42# a_n81_n130#
+ a_n321_n42# a_n509_n42# a_159_n42# a_351_n42# a_n33_n42# a_303_n130# a_n225_n42#
+ a_n177_64# a_207_64# a_n465_n130# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_n130# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_64# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n321_n42# a_n369_64# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n130# a_n509_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X8 a_n225_n42# a_n273_n130# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGLN5 a_n129_n130# a_n369_n42# a_1215_n130# a_543_64#
+ a_63_n130# a_159_64# a_n1089_n130# a_n849_n42# a_n417_64# a_n801_64# a_687_n42#
+ a_303_n42# a_1167_n42# a_n561_n42# a_n321_n130# a_n1041_n42# a_639_n130# a_n1185_64#
+ a_1023_n130# a_n1281_n130# a_n81_n42# a_399_n42# a_879_n42# a_n273_n42# a_735_64#
+ a_n753_n42# a_15_n42# a_n897_n130# a_n1233_n42# a_831_n130# a_447_n130# a_n609_64#
+ a_1071_n42# a_591_n42# a_1119_64# a_n993_64# a_207_n42# a_n465_n42# a_n945_n42#
+ a_351_64# a_783_n42# a_255_n130# a_n33_64# a_n225_64# a_n705_n130# a_1263_n42# a_927_64#
+ a_n177_n42# a_n657_n42# a_n1325_n42# a_n1137_n42# a_495_n42# a_111_n42# a_975_n42#
+ a_n513_n130# VSUBS
X0 a_303_n42# a_255_n130# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_591_n42# a_543_64# a_495_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_207_n42# a_159_64# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_399_n42# a_351_64# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_495_n42# a_447_n130# a_399_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_687_n42# a_639_n130# a_591_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_783_n42# a_735_64# a_687_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_975_n42# a_927_64# a_879_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n1041_n42# a_n1089_n130# a_n1137_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_879_n42# a_831_n130# a_783_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n1233_n42# a_n1281_n130# a_n1325_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X11 a_n1137_n42# a_n1185_64# a_n1233_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n561_n42# a_n609_64# a_n657_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1071_n42# a_1023_n130# a_975_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1263_n42# a_1215_n130# a_1167_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n945_n42# a_n993_64# a_n1041_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n753_n42# a_n801_64# a_n849_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n657_n42# a_n705_n130# a_n753_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n465_n42# a_n513_n130# a_n561_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n369_n42# a_n417_64# a_n465_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_1167_n42# a_1119_64# a_1071_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n849_n42# a_n897_n130# a_n945_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n273_n42# a_n321_n130# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n81_n42# a_n129_n130# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n177_n42# a_n225_64# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_VR4B8J a_1119_157# a_783_n126# a_n81_n126# a_n849_n126#
+ a_399_n126# a_n1041_n126# a_351_157# a_495_n126# a_n945_n126# a_n33_157# a_n129_n223#
+ a_n513_n223# a_1215_n223# a_63_n223# a_n1089_n223# a_n225_157# a_591_n126# a_n657_n126#
+ a_207_n126# a_543_157# a_n1325_n126# a_n369_n126# a_n753_n126# a_n321_n223# a_303_n126#
+ a_1023_n223# a_639_n223# a_n1281_n223# a_n417_157# a_n465_n126# a_1167_n126# a_735_157#
+ a_15_n126# a_n561_n126# a_n993_157# a_n177_n126# a_n897_n223# w_n1361_n226# a_1263_n126#
+ a_879_n126# a_111_n126# a_831_n223# a_n609_157# a_447_n223# a_n273_n126# a_n1137_n126#
+ a_975_n126# a_927_157# a_n1185_157# a_n1233_n126# a_n801_157# a_1071_n126# a_687_n126#
+ a_255_n223# a_n705_n223# a_159_157# VSUBS
X0 a_n273_n126# a_n321_n223# a_n369_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 a_n1233_n126# a_n1281_n223# a_n1325_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X2 a_591_n126# a_543_157# a_495_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 a_n849_n126# a_n897_n223# a_n945_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_207_n126# a_159_157# a_111_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_n177_n126# a_n225_157# a_n273_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X6 a_n1137_n126# a_n1185_157# a_n1233_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X7 a_495_n126# a_447_n223# a_399_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X8 a_n561_n126# a_n609_157# a_n657_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X9 a_111_n126# a_63_n223# a_15_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X10 a_783_n126# a_735_157# a_687_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X11 a_1071_n126# a_1023_n223# a_975_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X12 a_399_n126# a_351_157# a_303_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X13 a_n465_n126# a_n513_n223# a_n561_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X14 a_687_n126# a_639_n223# a_591_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X15 a_n753_n126# a_n801_157# a_n849_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X16 a_975_n126# a_927_157# a_879_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X17 a_n81_n126# a_n129_n223# a_n177_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X18 a_15_n126# a_n33_157# a_n81_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X19 a_1263_n126# a_1215_n223# a_1167_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X20 a_n1041_n126# a_n1089_n223# a_n1137_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X21 a_n369_n126# a_n417_157# a_n465_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X22 a_n657_n126# a_n705_n223# a_n753_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X23 a_879_n126# a_831_n223# a_783_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X24 a_n945_n126# a_n993_157# a_n1041_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X25 a_1167_n126# a_1119_157# a_1071_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X26 a_303_n126# a_255_n223# a_207_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
C0 w_n1361_n226# VSUBS 3.66914f
.ends

.subckt buffer a_1504_1398# m5_n1320_776# a_n1158_1778# a_1504_1860# a_1596_1398#
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS w_1358_2156# m4_n1330_2222#
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552#
+ a_n1158_1778# a_n1158_1778# a_1436_1552# a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_n1158_1778# a_1436_1552# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_1436_1552# a_1436_1552# a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552#
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_n1158_1778# a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# a_n1158_1778#
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_1436_1552# a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1778# w_1358_2156# a_1436_1552# a_1436_1552#
+ w_1358_2156# a_1436_1552# a_n1158_1778# a_1436_1552# w_1358_2156# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ w_1358_2156# a_1436_1552# w_1358_2156# a_n1158_1778# w_1358_2156# w_1358_2156# w_1358_2156#
+ a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ a_1436_1552# w_1358_2156# a_n1158_1778# w_1358_2156# w_1358_2156# a_n1158_1778#
+ w_1358_2156# a_n1158_1778# w_1358_2156# a_1436_1552# a_1436_1552# a_1436_1552# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_1436_1552# w_1358_2156# w_1358_2156# a_n1158_1778#
+ a_n1158_1778# a_1436_1552# a_n1158_1778# a_1436_1552# a_1436_1552# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
X0 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X2 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X6 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X8 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X11 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X12 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X15 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X16 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X17 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X20 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X21 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X24 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X27 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X30 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X32 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X35 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X36 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X38 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X39 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X43 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X45 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X46 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X48 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X49 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X50 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X53 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
C0 a_1596_1398# a_1504_1398# 2.6505f
C1 a_1504_1860# a_1596_1398# 6.786759f
C2 a_1436_1552# w_1358_2156# 4.344402f
C3 a_1436_1552# a_1596_1398# 2.21286f
C4 m5_n1320_776# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 2.587544f
C5 a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 8.208134f
C6 w_1358_2156# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 6.120336f
C7 a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 9.825851f
.ends

.subckt sky130_fd_pr__pfet_01v8_X4L24Q a_n33_n126# w_n353_n226# a_n317_n126# a_n177_157#
+ a_159_n126# a_111_n223# a_n273_n223# a_255_n126# a_n129_n126# a_n81_n223# a_63_n126#
+ a_n225_n126# a_15_157# a_207_157# VSUBS
X0 a_159_n126# a_111_n223# a_63_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 a_n225_n126# a_n273_n223# a_n317_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X2 a_63_n126# a_15_157# a_n33_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 a_n129_n126# a_n177_157# a_n225_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_n33_n126# a_n81_n223# a_n129_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_255_n126# a_207_157# a_159_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_XJUN3E a_63_n42# a_15_64# a_111_n130# a_n273_n130#
+ a_255_n42# a_n129_n42# a_n317_n42# a_n81_n130# a_159_n42# a_n33_n42# a_n225_n42#
+ a_n177_64# a_207_64# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n225_n42# a_n273_n130# a_n317_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X5 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt and_gate a_514_134# w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206#
+ m1_748_n50#
Xsky130_fd_pr__pfet_01v8_X4L24Q_0 w_n260_286# w_n260_286# m1_748_n50# a_n78_396# w_n260_286#
+ a_n78_396# a_n78_396# m1_748_n50# m1_748_n50# a_n78_396# m1_748_n50# w_n260_286#
+ a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q
Xsky130_fd_pr__nfet_01v8_XJUN3E_0 m1_748_n50# a_n78_396# a_n78_396# a_n78_396# m1_748_n50#
+ m1_748_n50# m1_748_n50# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__nfet_01v8_XJUN3E
X0 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.1953 pd=1.57 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_n78_396# a_514_134# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X6 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 w_n260_286# a_514_134# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.1953 ps=1.57 w=1.26 l=0.15
X8 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X9 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X10 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X11 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 w_n260_286# a_n78_396# 3.023118f
C1 a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 2.455001f
C2 w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 6.963798f
.ends

.subckt buffer_and_gate in1 clk out gnd vdd
Xbuffer_0 gnd gnd clk vdd m1_5444_838# gnd vdd vdd buffer
Xand_gate_0 m1_5444_838# vdd gnd in1 out and_gate
C0 in1 gnd 2.619732f
C1 and_gate_0/a_n78_396# gnd 2.338147f
C2 clk gnd 8.795321f
C3 m1_5444_838# gnd 2.352718f
C4 vdd gnd 18.256077f
C5 buffer_0/a_1436_1552# gnd 11.512064f
.ends

.subckt capacitor_5 cp_clk i1 vd2 vd1 vd4 vd3 clk GND VDD
Xbuffer_digital_1 i1 buffer_digital_1/in VDD GND buffer_digital_1/a_116_148# buffer_digital
Xsky130_fd_pr__nfet_01v8_D4CMYK_0 vd2 GND vd2 GND GND vd2 GND GND vd2 vd2 GND vd2
+ vd2 GND vd2 GND GND GND sky130_fd_pr__nfet_01v8_D4CMYK
Xsky130_fd_pr__pfet_01v8_4ZKXAA_1 vd3 vd3 GND vd3 vd3 GND vd3 GND vd3 GND GND vd3
+ GND vd3 vd3 GND GND vd3 vd3 GND vd3 GND GND sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__pfet_01v8_4ZKXAA_2 vd4 vd4 GND vd4 vd4 GND vd4 GND vd4 GND GND vd4
+ GND vd4 vd4 GND GND vd4 vd4 GND vd4 GND GND sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__pfet_01v8_4ZKXAA_3 vd3 vd3 GND vd3 vd3 GND vd3 GND vd3 GND GND vd3
+ GND vd3 vd3 GND GND vd3 vd3 GND vd3 GND GND sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__nfet_01v8_NJGC45_0 GND vd1 GND vd1 vd1 GND GND vd1 vd1 GND vd1 GND
+ GND GND GND GND vd1 GND vd1 vd1 vd1 GND sky130_fd_pr__nfet_01v8_NJGC45
Xbuffer_and_gate_0 buffer_digital_1/in clk buffer_and_gate_0/out GND VDD buffer_and_gate
X0 buffer_and_gate_0/out cp_clk sky130_fd_pr__cap_mim_m3_1 l=4.97 w=5
C0 i1 buffer_digital_1/in 2.935591f
C1 buffer_and_gate_0/and_gate_0/a_n78_396# GND 2.360761f
C2 clk GND 8.635434f
C3 VDD GND 20.988493f
C4 buffer_and_gate_0/buffer_0/a_1436_1552# GND 10.196393f
C5 vd1 GND 3.43263f
C6 vd3 GND 7.097779f
C7 vd4 GND 2.864619f
C8 vd2 GND 3.083021f
C9 buffer_digital_1/in GND 2.672912f
.ends

.subckt capacitors_5 capacitor_5_7/i1 capacitor_5_1/i1 capacitor_5_6/i1 capacitor_5_0/i1
+ capacitor_5_7/vd4 capacitor_5_3/i1 capacitor_5_7/vd2 capacitor_5_7/vd1 capacitor_5_7/cp_clk
+ capacitor_5_4/i1 capacitor_5_2/i1 capacitor_5_7/clk capacitor_5_7/vd3 capacitor_5_5/i1
+ capacitor_5_7/VDD VSUBS
Xcapacitor_5_5 capacitor_5_7/cp_clk capacitor_5_5/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_6 capacitor_5_7/cp_clk capacitor_5_6/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_7 capacitor_5_7/cp_clk capacitor_5_7/i1 capacitor_5_7/vd2 capacitor_5_7/vd1
+ capacitor_5_7/vd4 capacitor_5_7/vd3 capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_0 capacitor_5_7/cp_clk capacitor_5_0/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_1 capacitor_5_7/cp_clk capacitor_5_1/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_2 capacitor_5_7/cp_clk capacitor_5_2/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_3 capacitor_5_7/cp_clk capacitor_5_3/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_4 capacitor_5_7/cp_clk capacitor_5_4/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
C0 capacitor_5_7/VDD capacitor_5_7/clk 13.029696f
C1 capacitor_5_7/cp_clk capacitor_5_7/VDD 11.685536f
C2 capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.37575f
C3 capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.144792f
C4 capacitor_5_4/buffer_digital_1/in VSUBS 2.635156f
C5 capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.371064f
C6 capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.149221f
C7 capacitor_5_3/buffer_digital_1/in VSUBS 2.636791f
C8 capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.375672f
C9 capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.145726f
C10 capacitor_5_2/buffer_digital_1/in VSUBS 2.635774f
C11 capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.375235f
C12 capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.147629f
C13 capacitor_5_1/buffer_digital_1/in VSUBS 2.636666f
C14 capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C15 capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C16 capacitor_5_0/buffer_digital_1/in VSUBS 2.58165f
C17 capacitor_5_7/cp_clk VSUBS 20.068024f
C18 capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.376815f
C19 capacitor_5_7/clk VSUBS 71.174866f
C20 capacitor_5_7/VDD VSUBS 0.260321p
C21 capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.147582f
C22 capacitor_5_7/vd1 VSUBS 2.321869f
C23 capacitor_5_7/vd3 VSUBS 3.828029f
C24 capacitor_5_7/vd2 VSUBS 2.223177f
C25 capacitor_5_7/buffer_digital_1/in VSUBS 2.636351f
C26 capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.376023f
C27 capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.14572f
C28 capacitor_5_6/buffer_digital_1/in VSUBS 2.635363f
C29 capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.376738f
C30 capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.148531f
C31 capacitor_5_5/buffer_digital_1/in VSUBS 2.636503f
.ends

.subckt nmos_dnw3 vin out1 out2 clk clkb vs VSUBS
X0 clkb clk vin vs sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.126 ps=1.44 w=0.42 l=0.15
X1 vin clkb clk vs sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.1302 ps=1.46 w=0.42 l=0.15
X2 out2 clk vin vs sky130_fd_pr__nfet_01v8 ad=1.65 pd=7.1 as=0.945 ps=3.63 w=3 l=1
X3 vin clkb out1 vs sky130_fd_pr__nfet_01v8 ad=0.945 pd=3.63 as=1.65 ps=7.1 w=3 l=1
C0 vs VSUBS 6.63893f
.ends

.subckt sky130_fd_pr__pfet_01v8_FBZ64Q a_n81_n126# a_399_n126# a_351_n223# a_n417_n223#
+ a_207_n126# a_n225_n223# a_n461_n126# a_n369_n126# a_63_157# a_303_n126# a_255_157#
+ a_n33_n223# a_15_n126# a_n177_n126# a_n129_157# a_111_n126# w_n497_n226# a_n273_n126#
+ a_159_n223# a_n321_157# VSUBS
X0 a_n273_n126# a_n321_157# a_n369_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 a_207_n126# a_159_n223# a_111_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X2 a_n177_n126# a_n225_n223# a_n273_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 a_111_n126# a_63_157# a_15_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X4 a_399_n126# a_351_n223# a_303_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 a_n81_n126# a_n129_157# a_n177_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X6 a_15_n126# a_n33_n223# a_n81_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X7 a_n369_n126# a_n417_n223# a_n461_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X8 a_303_n126# a_255_157# a_207_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_5ACVEW a_n129_n130# a_63_n130# a_n81_n42# a_15_n42#
+ a_n173_n42# a_n33_64# a_111_n42# VSUBS
X0 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n81_n42# a_n129_n130# a_n173_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
.ends

.subckt inverter_27x m1_n804_1398# m1_540_1398# m1_156_1398# m1_n36_1398# m1_732_1398#
+ m1_n1102_1398# m1_348_1398# m1_n1188_1398# m1_n996_1398# m1_n228_1398# m1_n1188_1912#
+ m1_924_1398# m1_1309_1398# a_n1158_1658# m1_n420_1398# m1_1116_1398# w_1358_2036#
+ m1_n612_1398# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1658# m1_n228_1398# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# a_n1158_1658# a_n1158_1658#
+ m1_n1102_1398# m1_n1102_1398# m1_1309_1398# m1_n420_1398# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_540_1398#
+ m1_n1102_1398# m1_n1102_1398# a_n1158_1658# m1_n612_1398# m1_156_1398# a_n1158_1658#
+ m1_n1102_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_732_1398#
+ a_n1158_1658# a_n1158_1658# m1_348_1398# m1_n1102_1398# m1_n804_1398# a_n1158_1658#
+ m1_924_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# m1_n36_1398# m1_n1102_1398# m1_n1188_1398# m1_n996_1398# m1_n1102_1398#
+ m1_n1102_1398# m1_1116_1398# a_n1158_1658# VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1658# m1_n1188_1912# m1_1309_1398# m1_1309_1398#
+ m1_n1188_1912# m1_1309_1398# a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ m1_n1188_1912# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ a_n1158_1658# m1_n1188_1912# a_n1158_1658# w_1358_2036# m1_1309_1398# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_1309_1398# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# a_n1158_1658# m1_1309_1398# a_n1158_1658# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
C0 a_n1158_1658# VSUBS 6.394793f
C1 w_1358_2036# VSUBS 3.688076f
.ends

.subckt sky130_fd_pr__nfet_01v8_KMMFCM a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_29EZRJ a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_FL984Q a_n81_n126# a_n33_157# a_n129_n223# a_63_n223#
+ a_n173_n126# a_15_n126# a_111_n126# w_n209_n226# VSUBS
X0 a_111_n126# a_63_n223# a_15_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X1 a_n81_n126# a_n129_n223# a_n173_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X2 a_15_n126# a_n33_157# a_n81_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_D4CDWR a_n369_n42# a_n225_n130# a_303_n42# a_n81_n42#
+ a_399_n42# a_n33_n130# a_n273_n42# a_n461_n42# a_15_n42# a_n321_64# a_207_n42# a_159_n130#
+ a_n177_n42# a_351_n130# a_255_64# a_n417_n130# a_111_n42# a_n129_64# a_63_64# VSUBS
X0 a_303_n42# a_255_64# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_207_n42# a_159_n130# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_399_n42# a_351_n130# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n369_n42# a_n417_n130# a_n461_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X4 a_15_n42# a_n33_n130# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_111_n42# a_63_64# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n273_n42# a_n321_64# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n81_n42# a_n129_64# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n177_n42# a_n225_n130# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt clock clk_in vdd gnd clk clkb
Xsky130_fd_pr__pfet_01v8_FBZ64Q_0 vdd a_3246_118# a_2402_572# a_2402_572# a_3246_118#
+ a_2402_572# vdd a_3246_118# a_2402_572# vdd a_2402_572# a_2402_572# a_3246_118#
+ a_3246_118# a_2402_572# vdd vdd vdd a_2402_572# a_2402_572# gnd sky130_fd_pr__pfet_01v8_FBZ64Q
Xsky130_fd_pr__nfet_01v8_5ACVEW_0 a_344_n986# a_344_n986# a_2402_572# gnd gnd a_344_n986#
+ a_2402_572# gnd sky130_fd_pr__nfet_01v8_5ACVEW
Xinverter_27x_0 clk clk clk clk clk gnd clk clk clk clk vdd clk clk a_3246_118# clk
+ clk vdd clk gnd inverter_27x
Xsky130_fd_pr__nfet_01v8_KMMFCM_0 a_134_122# clk_in gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_1 a_416_120# a_344_102# sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42#
+ gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_2 sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42# a_134_122#
+ gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__pfet_01v8_29EZRJ_0 vdd vdd a_134_122# clk_in gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FL984Q_0 a_2402_572# a_344_n986# a_344_n986# a_344_n986#
+ vdd vdd a_2402_572# vdd gnd sky130_fd_pr__pfet_01v8_FL984Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 vdd vdd a_1230_122# m1_998_498# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_1 a_416_120# vdd vdd a_344_102# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 vdd vdd a_1430_122# a_1230_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_2 vdd vdd a_416_120# a_134_122# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_2 vdd vdd a_344_n986# a_1430_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_3 vdd vdd m1_998_498# a_786_n2# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__nfet_01v8_D4CDWR_0 a_3246_118# a_2402_572# gnd gnd a_3246_118# a_2402_572#
+ gnd gnd a_3246_118# a_2402_572# a_3246_118# a_2402_572# a_3246_118# a_2402_572#
+ a_2402_572# a_2402_572# gnd a_2402_572# a_2402_572# gnd sky130_fd_pr__nfet_01v8_D4CDWR
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 m1_998_498# a_786_n2# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 a_1230_122# m1_998_498# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_2 a_1430_122# a_1230_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_3 a_344_n986# a_1430_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
X0 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X2 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X3 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 vdd a_344_102# a_2020_n482# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X5 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X7 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X9 a_786_n912# a_586_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X10 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X11 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X12 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X13 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X17 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X20 a_286_n478# clk_in gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.15
X21 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X22 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X24 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_586_n2# a_416_120# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X27 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X28 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X30 a_786_n912# a_586_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X31 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X32 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 vdd a_344_n986# a_286_n960# vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.1827 ps=1.55 w=1.26 l=0.15
X34 a_344_102# a_1394_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X35 a_992_n918# a_786_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X36 a_1192_n918# a_992_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X37 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X38 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X39 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1394_n918# a_1192_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X42 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X43 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X46 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X48 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X49 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X51 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X52 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_586_n912# a_286_n960# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X54 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X55 a_586_n2# a_416_120# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X56 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X57 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X58 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X59 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X61 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X63 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X66 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X68 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_786_n2# a_586_n2# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X72 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_286_n960# clk_in vdd vdd sky130_fd_pr__pfet_01v8 ad=0.1827 pd=1.55 as=0.3654 ps=3.1 w=1.26 l=0.15
X74 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X75 a_286_n960# a_344_n986# a_286_n478# gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.15
X76 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X77 a_586_n912# a_286_n960# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X78 a_1394_n918# a_1192_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X79 a_1192_n918# a_992_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X80 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X81 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X82 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X83 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X84 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X85 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X86 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X87 a_344_102# a_1394_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X88 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.3906 ps=3.14 w=1.26 l=0.15
X89 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X90 gnd a_344_102# a_2020_n482# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X91 a_992_n918# a_786_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X92 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X93 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3906 pd=3.14 as=0.2079 ps=1.59 w=1.26 l=0.15
X94 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
X95 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X96 a_786_n2# a_586_n2# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X97 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.2079 pd=1.59 as=0.2079 ps=1.59 w=1.26 l=0.15
C0 a_2020_n482# vdd 2.656852f
C1 vdd clkb 7.306418f
C2 a_2432_n962# vdd 7.043292f
C3 a_2432_n962# clkb 2.67187f
C4 clkb gnd 5.097592f
C5 a_2432_n962# gnd 8.705547f
C6 a_2020_n482# gnd 2.565399f
C7 vdd gnd 26.103016f
C8 a_344_102# gnd 2.811321f
C9 a_2402_572# gnd 2.314155f
C10 a_344_n986# gnd 2.426004f
C11 a_3246_118# gnd 6.789812f
.ends

.subckt sky130_fd_pr__pfet_01v8_4RPJ49 a_2031_73# a_1887_n42# a_3615_n42# a_3183_73#
+ a_n3729_73# a_n2529_n42# a_1503_n42# a_63_n42# a_n753_n139# a_n3393_n42# a_n369_n139#
+ a_n1425_73# a_n1281_n42# a_n2961_73# a_687_73# a_n2577_73# a_n417_n42# a_2367_n42#
+ a_n1761_n42# a_n3009_n42# a_n2673_n139# a_2847_n42# a_n2289_n139# a_n3633_n139#
+ a_2607_73# a_n3249_n139# a_n1713_n139# a_3759_73# a_n1329_n139# a_255_n42# a_1455_73#
+ a_n2241_n42# a_2991_73# a_3471_n139# a_735_n42# a_1551_n139# a_3087_n139# a_1599_n42#
+ a_3327_n42# a_1167_n139# a_n2721_n42# a_n81_73# a_2511_n139# a_1215_n42# a_n273_73#
+ a_2127_n139# a_n993_n42# a_3807_n42# a_15_n139# a_303_73# a_n3585_n42# a_n129_n42#
+ a_2079_n42# a_n561_n139# a_n3345_73# a_n3201_n42# a_n1473_n42# a_n177_n139# a_n1041_73#
+ a_n609_n42# a_2559_n42# a_n2193_73# a_n1953_n42# a_n849_73# w_n3905_n142# a_n2481_n139#
+ a_n2097_n139# a_n3441_n139# a_1791_n42# a_n1521_n139# a_n3057_n139# a_2223_73# a_447_n42#
+ a_3039_n42# a_n1137_n139# a_3375_73# a_n2433_n42# a_927_n42# a_1071_73# a_n1617_73#
+ a_n2913_n42# a_3519_n42# a_975_n139# a_879_73# a_n2769_73# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n1185_n42# a_n801_n42# a_n3777_n42# a_2751_n42# a_n1665_n42#
+ a_1647_73# a_2799_73# a_3231_n42# a_159_n42# a_n2145_n42# a_n465_73# a_1983_n42#
+ a_3711_n42# a_639_n42# a_n2625_n42# a_1119_n42# a_n3537_73# a_n897_n42# a_n513_n42#
+ a_n1233_73# a_n3489_n42# a_2463_n42# a_783_n139# a_495_73# a_399_n139# a_n2385_73#
+ a_2895_n139# a_n3105_n42# a_n1377_n42# a_2943_n42# a_1935_n139# a_n1857_n42# a_351_n42#
+ a_2415_73# a_n33_n42# a_3567_73# a_831_n42# a_1695_n42# a_3423_n42# a_1263_73# a_n945_n139#
+ a_n2337_n42# a_1311_n42# a_n1809_73# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2175_n42#
+ a_n2865_n139# a_n1089_n42# a_n3825_n139# a_111_73# a_n2001_73# a_n3869_n42# a_n705_n42#
+ a_2655_n42# a_n1905_n139# a_n3153_73# a_591_n139# a_1839_73# a_n1569_n42# a_3663_n139#
+ a_1743_n139# a_3279_n139# a_543_n42# a_207_n139# a_n657_73# a_1359_n139# a_2703_n139#
+ a_3135_n42# VSUBS a_2319_n139# a_n2049_n42# a_1023_n42#
X0 a_n2241_n42# a_n2289_n139# a_n2337_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n2913_n42# a_n2961_73# a_n3009_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n2721_n42# a_n2769_73# a_n2817_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n2625_n42# a_n2673_n139# a_n2721_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n2433_n42# a_n2481_n139# a_n2529_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n2337_n42# a_n2385_73# a_n2433_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n2145_n42# a_n2193_73# a_n2241_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n2049_n42# a_n2097_n139# a_n2145_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n2817_n42# a_n2865_n139# a_n2913_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n2529_n42# a_n2577_73# a_n2625_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_2079_n42# a_2031_73# a_1983_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_2175_n42# a_2127_n139# a_2079_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_2271_n42# a_2223_73# a_2175_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_2367_n42# a_2319_n139# a_2271_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_2463_n42# a_2415_73# a_2367_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_2655_n42# a_2607_73# a_2559_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_2751_n42# a_2703_n139# a_2655_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_2943_n42# a_2895_n139# a_2847_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_2559_n42# a_2511_n139# a_2463_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_2847_n42# a_2799_73# a_2751_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_927_n42# a_879_73# a_831_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_1023_n42# a_975_n139# a_927_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n1953_n42# a_n2001_73# a_n2049_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_n1761_n42# a_n1809_73# a_n1857_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n1665_n42# a_n1713_n139# a_n1761_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n1857_n42# a_n1905_n139# a_n1953_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n1569_n42# a_n1617_73# a_n1665_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_1119_n42# a_1071_73# a_1023_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1215_n42# a_1167_n139# a_1119_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1311_n42# a_1263_73# a_1215_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_1407_n42# a_1359_n139# a_1311_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1503_n42# a_1455_73# a_1407_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_1695_n42# a_1647_73# a_1599_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1791_n42# a_1743_n139# a_1695_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1599_n42# a_1551_n139# a_1503_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_1887_n42# a_1839_73# a_1791_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_1983_n42# a_1935_n139# a_1887_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n33_n42# a_n81_73# a_n129_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_351_n42# a_303_73# a_255_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_159_n42# a_111_73# a_63_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_255_n42# a_207_n139# a_159_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_447_n42# a_399_n139# a_351_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_543_n42# a_495_73# a_447_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_639_n42# a_591_n139# a_543_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_735_n42# a_687_73# a_639_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_831_n42# a_783_n139# a_735_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_n1473_n42# a_n1521_n139# a_n1569_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_n1377_n42# a_n1425_73# a_n1473_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_n1281_n42# a_n1329_n139# a_n1377_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_n1185_n42# a_n1233_73# a_n1281_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n1089_n42# a_n1137_n139# a_n1185_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_n993_n42# a_n1041_73# a_n1089_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_n801_n42# a_n849_73# a_n897_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_n513_n42# a_n561_n139# a_n609_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_n321_n42# a_n369_n139# a_n417_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_n225_n42# a_n273_73# a_n321_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_n897_n42# a_n945_n139# a_n993_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_n705_n42# a_n753_n139# a_n801_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_n609_n42# a_n657_73# a_n705_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n417_n42# a_n465_73# a_n513_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n129_n42# a_n177_n139# a_n225_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_3327_n42# a_3279_n139# a_3231_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_3423_n42# a_3375_73# a_3327_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_3615_n42# a_3567_73# a_3519_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_3711_n42# a_3663_n139# a_3615_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_3519_n42# a_3471_n139# a_3423_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_3807_n42# a_3759_73# a_3711_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n3201_n42# a_n3249_n139# a_n3297_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_63_n42# a_15_n139# a_n33_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n3681_n42# a_n3729_73# a_n3777_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n3585_n42# a_n3633_n139# a_n3681_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n3393_n42# a_n3441_n139# a_n3489_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n3297_n42# a_n3345_73# a_n3393_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n3105_n42# a_n3153_73# a_n3201_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_n3009_n42# a_n3057_n139# a_n3105_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3231_n42# a_3183_73# a_3135_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_n3777_n42# a_n3825_n139# a_n3869_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X77 a_n3489_n42# a_n3537_73# a_n3585_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3039_n42# a_2991_73# a_2943_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3135_n42# a_3087_n139# a_3039_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 w_n3905_n142# VSUBS 6.63223f
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC8F a_15_n130# a_1887_n42# a_3615_n42# a_1647_64#
+ a_n561_n130# a_n2529_n42# a_1503_n42# a_2799_64# a_63_n42# a_n177_n130# a_n3393_n42#
+ a_n1281_n42# a_n465_64# a_n417_n42# a_2367_n42# a_n1761_n42# a_n2481_n130# a_n3009_n42#
+ a_n2097_n130# a_n3441_n130# a_2847_n42# a_n1521_n130# a_n3057_n130# a_n3537_64#
+ a_n1137_n130# a_255_n42# a_n1233_64# a_495_64# a_n2241_n42# a_n2385_64# a_975_n130#
+ a_735_n42# a_1599_n42# a_3327_n42# a_n2721_n42# a_1215_n42# a_2415_64# a_n993_n42#
+ a_3807_n42# a_3567_64# a_n3585_n42# a_n129_n42# a_2079_n42# a_1263_64# a_n3201_n42#
+ a_n1473_n42# a_n1809_64# a_n609_n42# a_2559_n42# a_n1953_n42# a_111_64# a_n2001_64#
+ a_1791_n42# a_447_n42# a_n3153_64# a_3039_n42# a_n2433_n42# a_1839_64# a_927_n42#
+ a_n2913_n42# a_3519_n42# a_783_n130# a_399_n130# a_2895_n130# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n657_64# a_n1185_n42# a_1935_n130# a_n801_n42# a_2031_64#
+ a_n3777_n42# a_2751_n42# a_3183_64# a_n1665_n42# a_n3729_64# a_n1425_64# a_687_64#
+ a_n2961_64# a_n945_n130# a_n2577_64# a_3231_n42# a_159_n42# a_n2145_n42# a_1983_n42#
+ a_3711_n42# a_2607_64# a_639_n42# a_n2625_n42# a_3759_64# a_n2865_n130# a_1119_n42#
+ a_n3825_n130# a_1455_64# a_n1905_n130# a_2991_64# a_n897_n42# a_591_n130# a_n513_n42#
+ a_n3489_n42# a_2463_n42# a_n3105_n42# a_n1377_n42# a_n81_64# a_n273_64# a_3663_n130#
+ a_3279_n130# a_2943_n42# a_1743_n130# a_207_n130# a_2703_n130# a_1359_n130# a_n1857_n42#
+ a_2319_n130# a_351_n42# a_303_64# a_n3345_64# a_n33_n42# a_831_n42# a_n1041_64#
+ a_1695_n42# a_3423_n42# a_n753_n130# a_n369_n130# a_n2193_64# a_n2337_n42# a_1311_n42#
+ a_n849_64# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2223_64# a_n2673_n130# a_2175_n42#
+ a_3375_64# a_n2289_n130# a_n3633_n130# a_n1089_n42# a_n3249_n130# a_n1713_n130#
+ a_n3869_n42# a_n705_n42# a_2655_n42# a_1071_64# a_n1329_n130# a_n1617_64# a_n1569_n42#
+ a_879_64# a_n2769_64# a_3471_n130# a_3087_n130# a_1551_n130# a_2511_n130# a_543_n42#
+ a_1167_n130# a_3135_n42# a_2127_n130# VSUBS a_n2049_n42# a_1023_n42#
X0 a_n3201_n42# a_n3249_n130# a_n3297_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n3681_n42# a_n3729_64# a_n3777_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n3585_n42# a_n3633_n130# a_n3681_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n3393_n42# a_n3441_n130# a_n3489_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n3297_n42# a_n3345_64# a_n3393_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n3105_n42# a_n3153_64# a_n3201_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n3009_n42# a_n3057_n130# a_n3105_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n3777_n42# a_n3825_n130# a_n3869_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X9 a_n3489_n42# a_n3537_64# a_n3585_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_3135_n42# a_3087_n130# a_3039_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_3231_n42# a_3183_64# a_3135_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_3039_n42# a_2991_64# a_2943_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n2241_n42# a_n2289_n130# a_n2337_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n2913_n42# a_n2961_64# a_n3009_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n2721_n42# a_n2769_64# a_n2817_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n2625_n42# a_n2673_n130# a_n2721_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n2433_n42# a_n2481_n130# a_n2529_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n2337_n42# a_n2385_64# a_n2433_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n2145_n42# a_n2193_64# a_n2241_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_n2049_n42# a_n2097_n130# a_n2145_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n2817_n42# a_n2865_n130# a_n2913_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n2529_n42# a_n2577_64# a_n2625_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2175_n42# a_2127_n130# a_2079_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_2271_n42# a_2223_64# a_2175_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2463_n42# a_2415_64# a_2367_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_2751_n42# a_2703_n130# a_2655_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_2079_n42# a_2031_64# a_1983_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_2367_n42# a_2319_n130# a_2271_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2559_n42# a_2511_n130# a_2463_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_2655_n42# a_2607_64# a_2559_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_2847_n42# a_2799_64# a_2751_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_2943_n42# a_2895_n130# a_2847_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1023_n42# a_975_n130# a_927_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_n1953_n42# a_n2001_64# a_n2049_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_n1761_n42# a_n1809_64# a_n1857_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n1665_n42# a_n1713_n130# a_n1761_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_n1857_n42# a_n1905_n130# a_n1953_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_n1569_n42# a_n1617_64# a_n1665_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1215_n42# a_1167_n130# a_1119_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1311_n42# a_1263_64# a_1215_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1503_n42# a_1455_64# a_1407_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_1791_n42# a_1743_n130# a_1695_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1119_n42# a_1071_64# a_1023_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_1407_n42# a_1359_n130# a_1311_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_1599_n42# a_1551_n130# a_1503_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1695_n42# a_1647_64# a_1599_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_1887_n42# a_1839_64# a_1791_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_1983_n42# a_1935_n130# a_1887_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n1473_n42# a_n1521_n130# a_n1569_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n1281_n42# a_n1329_n130# a_n1377_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_n1185_n42# a_n1233_64# a_n1281_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_n993_n42# a_n1041_64# a_n1089_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_n1377_n42# a_n1425_64# a_n1473_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_n1089_n42# a_n1137_n130# a_n1185_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n897_n42# a_n945_n130# a_n993_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_3327_n42# a_3279_n130# a_3231_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3423_n42# a_3375_64# a_3327_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_3615_n42# a_3567_64# a_3519_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X77 a_3711_n42# a_3663_n130# a_3615_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3519_n42# a_3471_n130# a_3423_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3807_n42# a_3759_64# a_3711_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt nmos_diode2 a_350_n764# a_970_n762# a_410_n892# dw_118_n1078# VSUBS
X0 a_410_n892# a_410_n892# a_350_n764# dw_118_n1078# sky130_fd_pr__nfet_01v8 ad=0.8729 pd=6.6 as=0.9029 ps=6.62 w=3.01 l=1
X1 a_350_n764# a_970_n762# a_970_n762# dw_118_n1078# sky130_fd_pr__nfet_01v8 ad=0.9929 pd=6.68 as=0.8729 ps=6.6 w=3.01 l=1
C0 dw_118_n1078# VSUBS 8.163819f
.ends

.subckt charge_pump in3 in5 input1 input2 out clk clkb clk_in g1 g2 vin in6 clock_0/vdd
+ in4 in8 in1 in7 clock_0/gnd in2 vs
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 g1 clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 g2 clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xcapacitors_5_1 in8 in2 in7 in1 clock_0/vdd in4 clock_0/vdd clock_0/vdd input2 in5
+ in3 clkb clock_0/vdd in6 clock_0/vdd clock_0/gnd capacitors_5
Xcapacitors_5_0 in8 in2 in7 in1 clock_0/vdd in4 clock_0/vdd clock_0/vdd input1 in5
+ in3 clk clock_0/vdd in6 clock_0/vdd clock_0/gnd capacitors_5
Xnmos_dnw3_0 vin input1 input2 g1 g2 vs clock_0/gnd nmos_dnw3
Xclock_0 clk_in clock_0/vdd clock_0/gnd clk clkb clock
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xnmos_diode2_0 out input2 input1 vs nmos_diode2_0/VSUBS nmos_diode2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 input2 clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 input1 clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 out clock_0/vdd 2.310455f
C1 vs input2 4.024266f
C2 vs clock_0/vdd 11.967723f
C3 vs clk 2.642354f
C4 clock_0/vdd clk 26.498407f
C5 vs input1 3.387235f
C6 input2 input1 8.763355f
C7 vs vin 8.809598f
C8 vs clkb 2.334149f
C9 vin clock_0/vdd 5.355844f
C10 clkb clock_0/vdd 17.402273f
C11 out vs 14.162664f
C12 vs nmos_diode2_0/VSUBS 20.067162f
C13 out nmos_diode2_0/VSUBS 3.142924f
C14 clock_0/a_2432_n962# nmos_diode2_0/VSUBS 8.684403f **FLOATING
C15 clock_0/a_2020_n482# nmos_diode2_0/VSUBS 2.571413f **FLOATING
C16 clock_0/a_344_102# nmos_diode2_0/VSUBS 2.810446f
C17 clock_0/a_2402_572# nmos_diode2_0/VSUBS 2.172722f
C18 clock_0/a_344_n986# nmos_diode2_0/VSUBS 2.381627f
C19 clock_0/a_3246_118# nmos_diode2_0/VSUBS 6.834443f
C20 g2 nmos_diode2_0/VSUBS 2.43748f
C21 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C22 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978447f
C23 capacitors_5_0/capacitor_5_4/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581751f
C24 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C25 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C26 capacitors_5_0/capacitor_5_3/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581653f
C27 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C28 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C29 capacitors_5_0/capacitor_5_2/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C30 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C31 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C32 capacitors_5_0/capacitor_5_1/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C33 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C34 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978566f
C35 capacitors_5_0/capacitor_5_0/buffer_digital_1/in nmos_diode2_0/VSUBS 2.583461f
C36 input1 nmos_diode2_0/VSUBS 16.681173f
C37 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C38 clk nmos_diode2_0/VSUBS 84.957054f
C39 clock_0/vdd nmos_diode2_0/VSUBS 0.459957p
C40 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978453f
C41 capacitors_5_0/capacitor_5_7/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581764f
C42 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C43 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978465f
C44 capacitors_5_0/capacitor_5_6/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581762f
C45 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C46 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978452f
C47 capacitors_5_0/capacitor_5_5/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581756f
C48 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C49 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C50 capacitors_5_1/capacitor_5_4/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C51 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C52 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.97846f
C53 capacitors_5_1/capacitor_5_3/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581745f
C54 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C55 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978502f
C56 capacitors_5_1/capacitor_5_2/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581764f
C57 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C58 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978491f
C59 capacitors_5_1/capacitor_5_1/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58176f
C60 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C61 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978744f
C62 capacitors_5_1/capacitor_5_0/buffer_digital_1/in nmos_diode2_0/VSUBS 2.583578f
C63 input2 nmos_diode2_0/VSUBS 16.89145f
C64 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C65 clkb nmos_diode2_0/VSUBS 87.08427f
C66 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C67 capacitors_5_1/capacitor_5_7/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581653f
C68 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C69 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C70 capacitors_5_1/capacitor_5_6/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C71 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.337696f
C72 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.978376f
C73 capacitors_5_1/capacitor_5_5/buffer_digital_1/in nmos_diode2_0/VSUBS 2.581652f
C74 g1 nmos_diode2_0/VSUBS 2.639545f
.ends

.subckt charge_pump_reverse m1_11946_n452# nmos_dnw3_0/out2 nmos_dnw3_0/vin clock_0/vdd
+ capacitors_5_1/capacitor_5_3/i1 clock_0/clk capacitors_5_1/capacitor_5_4/i1 clock_0/gnd
+ capacitors_5_1/capacitor_5_5/i1 capacitors_5_1/capacitor_5_2/i1 clock_0/clk_in capacitors_5_1/capacitor_5_7/i1
+ capacitors_5_1/capacitor_5_0/i1 capacitors_5_1/capacitor_5_6/i1 capacitors_5_1/capacitor_5_1/i1
+ nmos_dnw3_0/vs
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xcapacitors_5_1 capacitors_5_1/capacitor_5_7/i1 capacitors_5_1/capacitor_5_1/i1 capacitors_5_1/capacitor_5_6/i1
+ capacitors_5_1/capacitor_5_0/i1 clock_0/vdd capacitors_5_1/capacitor_5_3/i1 clock_0/vdd
+ clock_0/vdd nmos_dnw3_0/out2 capacitors_5_1/capacitor_5_4/i1 capacitors_5_1/capacitor_5_2/i1
+ clock_0/clk clock_0/vdd capacitors_5_1/capacitor_5_5/i1 clock_0/vdd clock_0/gnd
+ capacitors_5
Xcapacitors_5_0 capacitors_5_1/capacitor_5_7/i1 capacitors_5_1/capacitor_5_1/i1 capacitors_5_1/capacitor_5_6/i1
+ capacitors_5_1/capacitor_5_0/i1 clock_0/vdd capacitors_5_1/capacitor_5_3/i1 clock_0/vdd
+ clock_0/vdd nmos_dnw3_0/out1 capacitors_5_1/capacitor_5_4/i1 capacitors_5_1/capacitor_5_2/i1
+ clock_0/clkb clock_0/vdd capacitors_5_1/capacitor_5_5/i1 clock_0/vdd clock_0/gnd
+ capacitors_5
Xnmos_dnw3_0 nmos_dnw3_0/vin nmos_dnw3_0/out1 nmos_dnw3_0/out2 nmos_dnw3_0/clk nmos_dnw3_0/clkb
+ nmos_dnw3_0/vs clock_0/gnd nmos_dnw3
Xclock_0 clock_0/clk_in clock_0/vdd clock_0/gnd clock_0/clk clock_0/clkb clock
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xnmos_diode2_0 m1_11946_n452# nmos_dnw3_0/out2 nmos_dnw3_0/out1 nmos_dnw3_0/vs clock_0/gnd
+ nmos_diode2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 nmos_dnw3_0/out2 clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 nmos_dnw3_0/out1 clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 clock_0/vdd nmos_dnw3_0/vin 8.882092f
C1 clock_0/vdd clock_0/clk 20.03283f
C2 clock_0/vdd m1_11946_n452# 2.540002f
C3 clock_0/vdd nmos_dnw3_0/vs 2.471132f
C4 nmos_dnw3_0/out1 nmos_dnw3_0/out2 8.763353f
C5 m1_11946_n452# nmos_dnw3_0/vs 13.479089f
C6 nmos_dnw3_0/vs nmos_dnw3_0/out1 3.314235f
C7 nmos_dnw3_0/vs nmos_dnw3_0/out2 5.257541f
C8 clock_0/vdd clock_0/clkb 24.44572f
C9 nmos_dnw3_0/vs clock_0/gnd 19.463373f
C10 m1_11946_n452# clock_0/gnd 2.969539f
C11 clock_0/a_2432_n962# clock_0/gnd 8.689615f **FLOATING
C12 clock_0/a_2020_n482# clock_0/gnd 2.568188f **FLOATING
C13 clock_0/a_344_102# clock_0/gnd 2.809951f
C14 clock_0/a_2402_572# clock_0/gnd 2.172722f
C15 clock_0/a_344_n986# clock_0/gnd 2.381627f
C16 clock_0/a_3246_118# clock_0/gnd 6.834443f
C17 nmos_dnw3_0/vin clock_0/gnd 2.49859f
C18 nmos_dnw3_0/clkb clock_0/gnd 2.242713f
C19 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C20 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978447f
C21 capacitors_5_0/capacitor_5_4/buffer_digital_1/in clock_0/gnd 2.581751f
C22 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C23 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C24 capacitors_5_0/capacitor_5_3/buffer_digital_1/in clock_0/gnd 2.581652f
C25 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C26 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C27 capacitors_5_0/capacitor_5_2/buffer_digital_1/in clock_0/gnd 2.581652f
C28 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C29 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C30 capacitors_5_0/capacitor_5_1/buffer_digital_1/in clock_0/gnd 2.581652f
C31 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C32 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978566f
C33 capacitors_5_0/capacitor_5_0/buffer_digital_1/in clock_0/gnd 2.583461f
C34 nmos_dnw3_0/out1 clock_0/gnd 16.704819f
C35 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C36 clock_0/clkb clock_0/gnd 92.38439f
C37 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978453f
C38 capacitors_5_0/capacitor_5_7/buffer_digital_1/in clock_0/gnd 2.581764f
C39 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C40 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978465f
C41 capacitors_5_0/capacitor_5_6/buffer_digital_1/in clock_0/gnd 2.581762f
C42 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C43 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978452f
C44 capacitors_5_0/capacitor_5_5/buffer_digital_1/in clock_0/gnd 2.581756f
C45 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C46 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C47 capacitors_5_1/capacitor_5_4/buffer_digital_1/in clock_0/gnd 2.581652f
C48 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C49 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.97846f
C50 capacitors_5_1/capacitor_5_3/buffer_digital_1/in clock_0/gnd 2.581745f
C51 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C52 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978502f
C53 capacitors_5_1/capacitor_5_2/buffer_digital_1/in clock_0/gnd 2.581763f
C54 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C55 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978491f
C56 capacitors_5_1/capacitor_5_1/buffer_digital_1/in clock_0/gnd 2.58176f
C57 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C58 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978744f
C59 capacitors_5_1/capacitor_5_0/buffer_digital_1/in clock_0/gnd 2.583578f
C60 nmos_dnw3_0/out2 clock_0/gnd 16.02703f
C61 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C62 clock_0/clk clock_0/gnd 86.04303f
C63 clock_0/vdd clock_0/gnd 0.45817p
C64 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C65 capacitors_5_1/capacitor_5_7/buffer_digital_1/in clock_0/gnd 2.581653f
C66 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C67 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C68 capacitors_5_1/capacitor_5_6/buffer_digital_1/in clock_0/gnd 2.581652f
C69 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.337696f
C70 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.978376f
C71 capacitors_5_1/capacitor_5_5/buffer_digital_1/in clock_0/gnd 2.581652f
C72 nmos_dnw3_0/clk clock_0/gnd 2.52759f
.ends

.subckt CP2_5_stage charge_pump_reverse_1/nmos_dnw3_0/vs buffer_digital_7/in charge_pump_reverse_1/nmos_dnw3_0/out2
+ charge_pump_2/out charge_pump_0/out buffer_digital_7/VDD charge_pump_2/in3 charge_pump_0/vin
+ charge_pump_2/in4 charge_pump_reverse_1/clock_0/clk charge_pump_0/vs buffer_digital_4/i
+ charge_pump_2/in5 charge_pump_2/in6 charge_pump_1/vs charge_pump_reverse_0/nmos_dnw3_0/vs
+ charge_pump_2/in8 charge_pump_2/in1 buffer_digital_0/i buffer_digital_6/i buffer_digital_7/GND
+ charge_pump_2/in7 charge_pump_2/vs charge_pump_2/in2
Xcharge_pump_0 charge_pump_2/in3 charge_pump_2/in5 charge_pump_0/input1 charge_pump_0/input2
+ charge_pump_0/out charge_pump_0/clk charge_pump_0/clkb buffer_digital_0/i charge_pump_0/g1
+ charge_pump_0/g2 charge_pump_0/vin charge_pump_2/in6 buffer_digital_7/VDD charge_pump_2/in4
+ charge_pump_2/in8 charge_pump_2/in1 charge_pump_2/in7 buffer_digital_7/GND charge_pump_2/in2
+ charge_pump_0/vs charge_pump
Xcharge_pump_1 charge_pump_2/in3 charge_pump_2/in5 charge_pump_1/input1 charge_pump_1/input2
+ charge_pump_1/out charge_pump_1/clk charge_pump_1/clkb buffer_digital_4/i charge_pump_1/g1
+ charge_pump_1/g2 charge_pump_1/vin charge_pump_2/in6 buffer_digital_7/VDD charge_pump_2/in4
+ charge_pump_2/in8 charge_pump_2/in1 charge_pump_2/in7 buffer_digital_7/GND charge_pump_2/in2
+ charge_pump_1/vs charge_pump
Xbuffer_digital_0 buffer_digital_0/i buffer_digital_1/i buffer_digital_7/VDD buffer_digital_7/GND
+ buffer_digital_0/a_116_148# buffer_digital
Xcharge_pump_2 charge_pump_2/in3 charge_pump_2/in5 charge_pump_2/input1 charge_pump_2/input2
+ charge_pump_2/out charge_pump_2/clk charge_pump_2/clkb buffer_digital_7/in charge_pump_2/g1
+ charge_pump_2/g2 charge_pump_2/vin charge_pump_2/in6 buffer_digital_7/VDD charge_pump_2/in4
+ charge_pump_2/in8 charge_pump_2/in1 charge_pump_2/in7 buffer_digital_7/GND charge_pump_2/in2
+ charge_pump_2/vs charge_pump
Xbuffer_digital_1 buffer_digital_1/i buffer_digital_2/i buffer_digital_7/VDD buffer_digital_7/GND
+ buffer_digital_1/a_116_148# buffer_digital
Xbuffer_digital_2 buffer_digital_2/i buffer_digital_3/i buffer_digital_7/VDD buffer_digital_7/GND
+ buffer_digital_2/a_116_148# buffer_digital
Xbuffer_digital_3 buffer_digital_3/i buffer_digital_4/i buffer_digital_7/VDD buffer_digital_7/GND
+ buffer_digital_3/a_116_148# buffer_digital
Xbuffer_digital_5 buffer_digital_5/i buffer_digital_6/i buffer_digital_7/VDD buffer_digital_7/GND
+ buffer_digital_5/a_116_148# buffer_digital
Xbuffer_digital_4 buffer_digital_4/i buffer_digital_5/i buffer_digital_7/VDD buffer_digital_7/GND
+ buffer_digital_4/a_116_148# buffer_digital
Xbuffer_digital_6 buffer_digital_6/i buffer_digital_7/i buffer_digital_7/VDD buffer_digital_7/GND
+ buffer_digital_6/a_116_148# buffer_digital
Xbuffer_digital_7 buffer_digital_7/i buffer_digital_7/in buffer_digital_7/VDD buffer_digital_7/GND
+ buffer_digital_7/a_116_148# buffer_digital
Xcharge_pump_reverse_0 m2_44480_25420# charge_pump_reverse_0/nmos_dnw3_0/out2 charge_pump_0/out
+ buffer_digital_7/VDD charge_pump_2/in5 charge_pump_reverse_0/clock_0/clk charge_pump_2/in4
+ buffer_digital_7/GND charge_pump_2/in3 charge_pump_2/in6 buffer_digital_2/i charge_pump_2/in1
+ charge_pump_2/in8 charge_pump_2/in2 charge_pump_2/in7 charge_pump_reverse_0/nmos_dnw3_0/vs
+ charge_pump_reverse
Xcharge_pump_reverse_1 m2_91012_25410# charge_pump_reverse_1/nmos_dnw3_0/out2 charge_pump_1/out
+ buffer_digital_7/VDD charge_pump_2/in5 charge_pump_reverse_1/clock_0/clk charge_pump_2/in4
+ buffer_digital_7/GND charge_pump_2/in3 charge_pump_2/in6 buffer_digital_6/i charge_pump_2/in1
+ charge_pump_2/in8 charge_pump_2/in2 charge_pump_2/in7 charge_pump_reverse_1/nmos_dnw3_0/vs
+ charge_pump_reverse
C0 buffer_digital_7/VDD buffer_digital_4/i 4.262721f
C1 buffer_digital_7/VDD charge_pump_2/in2 4.191784f
C2 buffer_digital_7/VDD charge_pump_2/in5 4.276729f
C3 buffer_digital_7/VDD charge_pump_2/in7 4.29743f
C4 buffer_digital_7/VDD buffer_digital_6/i 4.442357f
C5 buffer_digital_7/VDD charge_pump_2/in4 4.281688f
C6 buffer_digital_7/VDD charge_pump_2/in1 4.123556f
C7 buffer_digital_7/VDD charge_pump_2/in6 4.186176f
C8 buffer_digital_7/VDD buffer_digital_7/in 2.184147f
C9 buffer_digital_7/VDD charge_pump_2/in3 4.304672f
C10 buffer_digital_7/VDD buffer_digital_2/i 4.399636f
C11 buffer_digital_7/VDD charge_pump_2/in8 4.333586f
C12 buffer_digital_7/VDD buffer_digital_0/i 4.540237f
C13 charge_pump_reverse_1/nmos_dnw3_0/vs buffer_digital_7/GND 18.799433f
C14 charge_pump_reverse_1/clock_0/a_2432_n962# buffer_digital_7/GND 8.68424f **FLOATING
C15 charge_pump_reverse_1/clock_0/a_2020_n482# buffer_digital_7/GND 2.56615f **FLOATING
C16 charge_pump_reverse_1/clock_0/a_344_102# buffer_digital_7/GND 2.809951f
C17 charge_pump_reverse_1/clock_0/a_2402_572# buffer_digital_7/GND 2.172722f
C18 charge_pump_reverse_1/clock_0/a_344_n986# buffer_digital_7/GND 2.381627f
C19 charge_pump_reverse_1/clock_0/a_3246_118# buffer_digital_7/GND 6.834443f
C20 charge_pump_reverse_1/nmos_dnw3_0/clkb buffer_digital_7/GND 2.234749f
C21 charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C22 charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C23 charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C24 charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C25 charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C26 charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C27 charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C28 charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C29 charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C30 charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C31 charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C32 charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C33 charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C34 charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C35 charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C36 charge_pump_reverse_1/nmos_dnw3_0/out1 buffer_digital_7/GND 15.064581f
C37 charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C38 charge_pump_reverse_1/clock_0/clkb buffer_digital_7/GND 91.19051f
C39 charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C40 charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C41 charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C42 charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C43 charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C44 charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C45 charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C46 charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C47 charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C48 charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C49 charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C50 charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C51 charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C52 charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C53 charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C54 charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C55 charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C56 charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C57 charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C58 charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C59 charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C60 charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C61 charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C62 charge_pump_reverse_1/nmos_dnw3_0/out2 buffer_digital_7/GND 14.843945f
C63 charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C64 charge_pump_reverse_1/clock_0/clk buffer_digital_7/GND 84.467705f
C65 charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C66 charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C67 charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C68 charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C69 charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C70 charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C71 charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C72 charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C73 charge_pump_reverse_1/nmos_dnw3_0/clk buffer_digital_7/GND 2.425359f
C74 charge_pump_reverse_0/nmos_dnw3_0/vs buffer_digital_7/GND 18.80054f
C75 charge_pump_reverse_0/clock_0/a_2432_n962# buffer_digital_7/GND 8.68424f **FLOATING
C76 charge_pump_reverse_0/clock_0/a_2020_n482# buffer_digital_7/GND 2.56615f **FLOATING
C77 charge_pump_reverse_0/clock_0/a_344_102# buffer_digital_7/GND 2.809951f
C78 charge_pump_reverse_0/clock_0/a_2402_572# buffer_digital_7/GND 2.172722f
C79 charge_pump_reverse_0/clock_0/a_344_n986# buffer_digital_7/GND 2.381627f
C80 charge_pump_reverse_0/clock_0/a_3246_118# buffer_digital_7/GND 6.834443f
C81 charge_pump_reverse_0/nmos_dnw3_0/clkb buffer_digital_7/GND 2.234749f
C82 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C83 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C84 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C85 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C86 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C87 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C88 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C89 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C90 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C91 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C92 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C93 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C94 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C95 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C96 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C97 charge_pump_reverse_0/nmos_dnw3_0/out1 buffer_digital_7/GND 15.064581f
C98 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C99 charge_pump_reverse_0/clock_0/clkb buffer_digital_7/GND 91.13845f
C100 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C101 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C102 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C103 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C104 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C105 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C106 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C107 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C108 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C109 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C110 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C111 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C112 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C113 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C114 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C115 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C116 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C117 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C118 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C119 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C120 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C121 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C122 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C123 charge_pump_reverse_0/nmos_dnw3_0/out2 buffer_digital_7/GND 14.843945f
C124 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C125 charge_pump_reverse_0/clock_0/clk buffer_digital_7/GND 84.59574f
C126 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C127 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C128 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C129 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C130 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C131 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C132 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C133 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C134 charge_pump_reverse_0/nmos_dnw3_0/clk buffer_digital_7/GND 2.425359f
C135 buffer_digital_6/i buffer_digital_7/GND 10.521893f
C136 buffer_digital_2/i buffer_digital_7/GND 8.909059f
C137 charge_pump_2/vs buffer_digital_7/GND 18.96316f
C138 charge_pump_2/clock_0/a_2432_n962# buffer_digital_7/GND 8.68424f **FLOATING
C139 charge_pump_2/clock_0/a_2020_n482# buffer_digital_7/GND 2.56615f **FLOATING
C140 charge_pump_2/clock_0/a_344_102# buffer_digital_7/GND 2.809951f
C141 charge_pump_2/clock_0/a_2402_572# buffer_digital_7/GND 2.172722f
C142 charge_pump_2/clock_0/a_344_n986# buffer_digital_7/GND 2.381627f
C143 buffer_digital_7/in buffer_digital_7/GND 17.948488f
C144 charge_pump_2/clock_0/a_3246_118# buffer_digital_7/GND 6.834443f
C145 charge_pump_2/g2 buffer_digital_7/GND 2.43748f
C146 charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C147 charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C148 charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C149 charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C150 charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C151 charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C152 charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C153 charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C154 charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C155 charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C156 charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C157 charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C158 charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C159 charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C160 charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C161 charge_pump_2/in1 buffer_digital_7/GND 13.808674f
C162 charge_pump_2/input1 buffer_digital_7/GND 15.031953f
C163 charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C164 charge_pump_2/clk buffer_digital_7/GND 82.25474f
C165 charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C166 charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C167 charge_pump_2/in8 buffer_digital_7/GND 13.756854f
C168 charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C169 charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C170 charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C171 charge_pump_2/in7 buffer_digital_7/GND 14.582843f
C172 charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C173 charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C174 charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C175 charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C176 charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C177 charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C178 charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C179 charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C180 charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C181 charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C182 charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C183 charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C184 charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C185 charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C186 charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C187 charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C188 charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C189 charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C190 charge_pump_2/input2 buffer_digital_7/GND 14.390842f
C191 charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C192 charge_pump_2/clkb buffer_digital_7/GND 83.97966f
C193 charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C194 charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C195 charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C196 charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C197 charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C198 charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C199 charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C200 charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C201 charge_pump_2/g1 buffer_digital_7/GND 2.634558f
C202 buffer_digital_1/i buffer_digital_7/GND 2.411286f
C203 charge_pump_1/vs buffer_digital_7/GND 18.977581f
C204 charge_pump_1/out buffer_digital_7/GND 3.739746f
C205 charge_pump_1/clock_0/a_2432_n962# buffer_digital_7/GND 8.68424f **FLOATING
C206 charge_pump_1/clock_0/a_2020_n482# buffer_digital_7/GND 2.56615f **FLOATING
C207 charge_pump_1/clock_0/a_344_102# buffer_digital_7/GND 2.809951f
C208 charge_pump_1/clock_0/a_2402_572# buffer_digital_7/GND 2.172722f
C209 charge_pump_1/clock_0/a_344_n986# buffer_digital_7/GND 2.381627f
C210 buffer_digital_4/i buffer_digital_7/GND 14.695759f
C211 charge_pump_1/clock_0/a_3246_118# buffer_digital_7/GND 6.834443f
C212 charge_pump_1/g2 buffer_digital_7/GND 2.43748f
C213 charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C214 charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C215 charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C216 charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C217 charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C218 charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C219 charge_pump_2/in4 buffer_digital_7/GND 14.559189f
C220 charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C221 charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C222 charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C223 charge_pump_2/in3 buffer_digital_7/GND 14.574407f
C224 charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C225 charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C226 charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C227 charge_pump_2/in2 buffer_digital_7/GND 14.538905f
C228 charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C229 charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C230 charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C231 charge_pump_1/input1 buffer_digital_7/GND 15.031953f
C232 charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C233 charge_pump_1/clk buffer_digital_7/GND 82.53111f
C234 charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C235 charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C236 charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C237 charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C238 charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C239 charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C240 charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C241 charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C242 charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C243 charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C244 charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C245 charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C246 charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C247 charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C248 charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C249 charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C250 charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C251 charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C252 charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C253 charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C254 charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C255 charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C256 charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C257 charge_pump_1/input2 buffer_digital_7/GND 14.390842f
C258 charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C259 charge_pump_1/clkb buffer_digital_7/GND 84.08535f
C260 charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C261 charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C262 charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C263 charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C264 charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C265 charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C266 charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C267 charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C268 charge_pump_1/g1 buffer_digital_7/GND 2.634558f
C269 charge_pump_0/vs buffer_digital_7/GND 18.974451f
C270 charge_pump_0/out buffer_digital_7/GND 2.335674f
C271 charge_pump_0/clock_0/a_2432_n962# buffer_digital_7/GND 8.68424f **FLOATING
C272 charge_pump_0/clock_0/a_2020_n482# buffer_digital_7/GND 2.56615f **FLOATING
C273 charge_pump_0/clock_0/a_344_102# buffer_digital_7/GND 2.809951f
C274 charge_pump_0/clock_0/a_2402_572# buffer_digital_7/GND 2.172722f
C275 charge_pump_0/clock_0/a_344_n986# buffer_digital_7/GND 2.381627f
C276 buffer_digital_0/i buffer_digital_7/GND 17.110367f
C277 charge_pump_0/clock_0/a_3246_118# buffer_digital_7/GND 6.834443f
C278 charge_pump_0/g2 buffer_digital_7/GND 2.43748f
C279 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C280 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C281 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C282 charge_pump_2/in5 buffer_digital_7/GND 14.567261f
C283 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C284 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C285 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C286 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C287 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C288 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C289 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C290 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C291 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C292 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C293 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C294 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C295 charge_pump_0/input1 buffer_digital_7/GND 15.031953f
C296 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C297 charge_pump_0/clk buffer_digital_7/GND 82.54194f
C298 buffer_digital_7/VDD buffer_digital_7/GND 2.225115p
C299 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C300 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C301 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C302 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C303 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C304 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C305 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C306 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C307 charge_pump_2/in6 buffer_digital_7/GND 14.385935f
C308 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C309 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C310 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C311 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C312 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C313 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C314 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C315 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C316 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C317 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C318 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C319 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C320 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C321 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C322 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C323 charge_pump_0/input2 buffer_digital_7/GND 14.391004f
C324 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C325 charge_pump_0/clkb buffer_digital_7/GND 84.04496f
C326 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C327 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C328 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C329 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C330 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C331 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# buffer_digital_7/GND 2.337696f
C332 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# buffer_digital_7/GND 9.978376f
C333 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in buffer_digital_7/GND 2.581652f
C334 charge_pump_0/g1 buffer_digital_7/GND 2.634558f
.ends

.subckt sky130_fd_pr__nfet_01v8_9LGCGE a_15_n130# a_n561_n130# a_63_n42# a_n989_n42#
+ a_n177_n130# a_n417_n42# a_n465_64# a_255_n42# a_495_64# a_735_n42# a_n129_n42#
+ a_n609_n42# a_111_64# a_447_n42# a_927_n42# a_783_n130# a_n321_n42# a_399_n130#
+ a_n657_64# a_n801_n42# a_687_64# a_n945_n130# a_159_n42# a_639_n42# a_n513_n42#
+ a_n897_n42# a_591_n130# a_n81_64# a_n273_64# a_351_n42# a_207_n130# a_303_64# a_n33_n42#
+ a_831_n42# a_n369_n130# a_n753_n130# a_n849_64# a_n225_n42# a_n705_n42# a_879_64#
+ a_543_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n897_n42# a_n945_n130# a_n989_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_49FP49 a_63_n42# a_n989_n42# a_n369_n139# a_n753_n139#
+ a_n417_n42# a_687_73# w_n1025_n142# a_255_n42# a_735_n42# a_n81_73# a_n273_73# a_n129_n42#
+ a_15_n139# a_n561_n139# a_303_73# a_n609_n42# a_n177_n139# a_n849_73# a_447_n42#
+ a_927_n42# a_n321_n42# a_879_73# a_n801_n42# a_159_n42# a_639_n42# a_n465_73# a_n513_n42#
+ a_n897_n42# a_783_n139# a_495_73# a_399_n139# a_351_n42# a_n33_n42# a_831_n42# a_n945_n139#
+ a_n225_n42# a_n705_n42# a_111_73# a_591_n139# a_543_n42# a_207_n139# a_n657_73#
+ VSUBS
X0 a_927_n42# a_879_73# a_831_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_73# a_n129_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_73# a_255_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_73# a_63_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n139# a_159_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_n139# a_351_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_543_n42# a_495_73# a_447_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_639_n42# a_591_n139# a_543_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_73# a_639_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n139# a_735_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n801_n42# a_n849_73# a_n897_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n513_n42# a_n561_n139# a_n609_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n321_n42# a_n369_n139# a_n417_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n225_n42# a_n273_73# a_n321_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n897_n42# a_n945_n139# a_n989_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X15 a_n705_n42# a_n753_n139# a_n801_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n609_n42# a_n657_73# a_n705_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n417_n42# a_n465_73# a_n513_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n139# a_n225_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_63_n42# a_15_n139# a_n33_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt capacito7 a_2858_n174# sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142# buffer_digital_0/i
+ a_5270_n124# m3_7758_166# buffer_and_gate_0/clk sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142#
+ m1_6370_n278# buffer_digital_0/VDD m1_602_n334# VSUBS
Xbuffer_digital_0 buffer_digital_0/i buffer_digital_0/in buffer_digital_0/VDD VSUBS
+ buffer_digital_0/a_116_148# buffer_digital
Xsky130_fd_pr__pfet_01v8_4ZKXAA_0 m1_6370_n278# m1_6370_n278# VSUBS sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142#
+ m1_6370_n278# VSUBS m1_6370_n278# VSUBS m1_6370_n278# VSUBS VSUBS m1_6370_n278#
+ VSUBS m1_6370_n278# m1_6370_n278# VSUBS VSUBS m1_6370_n278# m1_6370_n278# VSUBS
+ m1_6370_n278# VSUBS VSUBS sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__nfet_01v8_9LGCGE_0 a_2858_n174# a_2858_n174# VSUBS VSUBS a_2858_n174#
+ VSUBS a_2858_n174# VSUBS a_2858_n174# VSUBS VSUBS VSUBS a_2858_n174# VSUBS VSUBS
+ a_2858_n174# VSUBS a_2858_n174# a_2858_n174# VSUBS a_2858_n174# a_2858_n174# VSUBS
+ VSUBS VSUBS VSUBS a_2858_n174# a_2858_n174# a_2858_n174# VSUBS a_2858_n174# a_2858_n174#
+ VSUBS VSUBS a_2858_n174# a_2858_n174# a_2858_n174# VSUBS VSUBS a_2858_n174# VSUBS
+ VSUBS sky130_fd_pr__nfet_01v8_9LGCGE
Xsky130_fd_pr__pfet_01v8_49FP49_0 m1_602_n334# m1_602_n334# VSUBS VSUBS m1_602_n334#
+ VSUBS sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142# m1_602_n334# m1_602_n334# VSUBS
+ VSUBS m1_602_n334# VSUBS VSUBS VSUBS m1_602_n334# VSUBS VSUBS m1_602_n334# m1_602_n334#
+ m1_602_n334# VSUBS m1_602_n334# m1_602_n334# m1_602_n334# VSUBS m1_602_n334# m1_602_n334#
+ VSUBS VSUBS VSUBS m1_602_n334# m1_602_n334# m1_602_n334# VSUBS m1_602_n334# m1_602_n334#
+ VSUBS VSUBS m1_602_n334# VSUBS VSUBS VSUBS sky130_fd_pr__pfet_01v8_49FP49
Xsky130_fd_pr__nfet_01v8_NJGC45_0 VSUBS a_5270_n124# VSUBS a_5270_n124# a_5270_n124#
+ VSUBS VSUBS a_5270_n124# a_5270_n124# VSUBS a_5270_n124# VSUBS VSUBS VSUBS VSUBS
+ VSUBS a_5270_n124# VSUBS a_5270_n124# a_5270_n124# a_5270_n124# VSUBS sky130_fd_pr__nfet_01v8_NJGC45
Xbuffer_and_gate_0 buffer_digital_0/in buffer_and_gate_0/clk buffer_and_gate_0/out
+ VSUBS buffer_digital_0/VDD buffer_and_gate
X0 buffer_and_gate_0/out m3_7758_166# sky130_fd_pr__cap_mim_m3_1 l=7.99 w=7.97
C0 buffer_digital_0/in buffer_digital_0/i 2.942645f
C1 m3_7758_166# VSUBS 2.50035f
C2 buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.473223f
C3 buffer_and_gate_0/clk VSUBS 8.924417f
C4 buffer_digital_0/VDD VSUBS 18.041912f
C5 buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.15507f
C6 a_5270_n124# VSUBS 3.420046f
C7 m1_602_n334# VSUBS 2.778242f
C8 a_2858_n174# VSUBS 6.69811f
C9 buffer_digital_0/in VSUBS 2.681842f
.ends

.subckt capacitor_8 capacitor_7_0/a_5270_n124# capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/clk
+ capacitor_7_0/buffer_digital_0/VDD capacitor_7_0/a_2858_n174# w_7118_n356# w_1380_n364#
+ VSUBS capacitor_7_0/buffer_digital_0/i
Xcapacitor_7_0 capacitor_7_0/a_2858_n174# w_7118_n356# capacitor_7_0/buffer_digital_0/i
+ capacitor_7_0/a_5270_n124# capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/clk
+ w_1380_n364# w_7118_n356# capacitor_7_0/buffer_digital_0/VDD w_1380_n364# VSUBS
+ capacito7
C0 capacitor_7_0/m3_7758_166# VSUBS 2.31534f
C1 capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C2 capacitor_7_0/buffer_and_gate_0/clk VSUBS 8.196827f
C3 capacitor_7_0/buffer_digital_0/VDD VSUBS 18.215277f
C4 capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C5 capacitor_7_0/a_5270_n124# VSUBS 2.356963f
C6 w_1380_n364# VSUBS 3.53509f
C7 capacitor_7_0/a_2858_n174# VSUBS 4.668162f
C8 capacitor_7_0/buffer_digital_0/in VSUBS 2.608221f
.ends

.subckt capacitors_1 clk1 capacitor_8_0/capacitor_7_0/a_2858_n174# capacitor_8_0/capacitor_7_0/a_5270_n124#
+ capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk capacitor_8_0/capacitor_7_0/buffer_digital_0/VDD
+ m1_7096_n308# capacitor_8_0/w_1380_n364# in1 VSUBS
Xcapacitor_8_0 capacitor_8_0/capacitor_7_0/a_5270_n124# clk1 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk
+ capacitor_8_0/capacitor_7_0/buffer_digital_0/VDD capacitor_8_0/capacitor_7_0/a_2858_n174#
+ m1_7096_n308# capacitor_8_0/w_1380_n364# VSUBS in1 capacitor_8
C0 clk1 VSUBS 2.376945f
C1 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.337696f
C2 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk VSUBS 9.493001f
C3 capacitor_8_0/capacitor_7_0/buffer_digital_0/VDD VSUBS 22.92377f
C4 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.978376f
C5 capacitor_8_0/capacitor_7_0/a_5270_n124# VSUBS 2.356963f
C6 capacitor_8_0/w_1380_n364# VSUBS 3.265198f
C7 capacitor_8_0/capacitor_7_0/a_2858_n174# VSUBS 4.668162f
C8 capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.613958f
.ends

.subckt sky130_fd_pr__pfet_01v8_E9H44Q a_15_n42# a_n15_n68# w_n109_n104# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# w_n109_n104# sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_9AYYDL a_n158_n300# w_n194_n362# a_100_n300# a_n100_n326#
+ VSUBS
X0 a_100_n300# a_n100_n326# a_n158_n300# w_n194_n362# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt pmos_cp1 a_168_22# m1_532_58# w_n14_n142# a_424_18# m1_14_56# VSUBS
Xsky130_fd_pr__pfet_01v8_E9H44Q_0 w_n14_n142# a_168_22# w_n14_n142# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_E9H44Q_1 a_168_22# a_424_18# w_n14_n142# w_n14_n142# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_9AYYDL_0 m1_14_56# w_n14_n142# w_n14_n142# a_168_22# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
Xsky130_fd_pr__pfet_01v8_9AYYDL_1 w_n14_n142# w_n14_n142# m1_532_58# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
C0 w_n14_n142# VSUBS 2.470929f
.ends

.subckt charge_pump1 clk_in input1 input2 vdd in1 in2 in6 in7 g1 g2 clk clkb m1_12464_n576#
+ a_3340_18086# in4 gnd in3 in5 in8 vin
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 g1 clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 g2 clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 vin input1 input2 g1 g2 vin gnd nmos_dnw3
Xclock_0 clk_in vdd gnd clk clkb clock
Xcapacitor_8_0 vdd input1 clk vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 clkb vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 vdd vdd clk vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_1 input2 vdd vdd clkb vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_2 input1 vdd vdd clk vdd vdd vdd in2 gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 vdd vdd clk vdd vdd vdd in3 gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_4 input2 vdd vdd clkb vdd vdd vdd in2 gnd capacitors_1
Xcapacitors_1_5 input2 vdd vdd clkb vdd vdd vdd in3 gnd capacitors_1
Xcapacitors_1_6 input1 vdd vdd clk vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_7 input1 vdd vdd clk vdd vdd vdd in5 gnd capacitors_1
Xcapacitors_1_8 input1 vdd vdd clk vdd vdd vdd in6 gnd capacitors_1
Xcapacitors_1_9 input1 vdd vdd clk vdd vdd vdd in7 gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 vdd vdd clkb vdd vdd vdd in7 gnd capacitors_1
Xcapacitors_1_11 input2 vdd vdd clkb vdd vdd vdd in6 gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 vdd vdd clkb vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_12 input2 vdd vdd clkb vdd vdd vdd in5 gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clkb input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clk input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 clk m1_12464_n576# 2.312213f
C1 clkb m1_12464_n576# 2.207061f
C2 input2 vdd 26.500193f
C3 vdd vin 9.1372f
C4 vin clk 2.188878f
C5 input2 input1 3.059187f
C6 vdd clk 32.205326f
C7 input1 vdd 26.823656f
C8 vdd clkb 26.212053f
C9 input1 gnd 30.964584f
C10 input2 gnd 31.05456f
C11 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.396566f
C12 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.07966f
C13 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634299f
C14 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398093f
C15 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.08029f
C16 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633591f
C17 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.392522f
C18 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079402f
C19 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634253f
C20 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398324f
C21 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079739f
C22 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633955f
C23 m1_4341_n519# gnd 4.097057f
C24 m1_12659_300# gnd 2.789905f
C25 m1_12464_n576# gnd 5.227879f
C26 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.397358f
C27 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079556f
C28 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634405f
C29 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.394424f
C30 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079654f
C31 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634067f
C32 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393486f
C33 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.07973f
C34 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633915f
C35 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393389f
C36 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079822f
C37 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633871f
C38 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398049f
C39 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079473f
C40 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633938f
C41 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.396035f
C42 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079795f
C43 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634021f
C44 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.395022f
C45 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079731f
C46 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634052f
C47 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.392135f
C48 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.078752f
C49 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633513f
C50 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.338151f
C51 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.97841f
C52 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61055f
C53 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.33782f
C54 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978384f
C55 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.610197f
C56 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393725f
C57 clkb gnd 91.86899f
C58 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.080707f
C59 capacitor_8_1/capacitor_7_0/buffer_digital_0/in gnd 2.639488f
C60 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.397516f
C61 clk gnd 91.63095f
C62 vdd gnd 0.653035p
C63 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079217f
C64 capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.639593f
C65 clock_0/a_2432_n962# gnd 8.68424f **FLOATING
C66 clock_0/a_2020_n482# gnd 2.567662f **FLOATING
C67 clock_0/a_344_102# gnd 2.813001f
C68 clock_0/a_2402_572# gnd 2.172722f
C69 clock_0/a_344_n986# gnd 2.381627f
C70 clock_0/a_3246_118# gnd 6.834443f
C71 g2 gnd 2.344427f
C72 vin gnd 10.416249f
.ends

.subckt charge_pump1_reverse input1 input2 in1 in2 in6 in7 vdd m1_12464_n576# clock_1/clk_in
+ a_3340_18086# gnd in4 in3 in5 in8 nmos_dnw3_0/vs
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 nmos_dnw3_0/vs input1 input2 nmos_dnw3_0/clk nmos_dnw3_0/clkb nmos_dnw3_0/vs
+ gnd nmos_dnw3
Xclock_1 clock_1/clk_in vdd gnd clock_1/clk clock_1/clkb clock
Xcapacitor_8_0 vdd input1 clock_1/clkb vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 clock_1/clk vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 vdd vdd clock_1/clkb vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_1 input2 vdd vdd clock_1/clk vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_2 input1 vdd vdd clock_1/clkb vdd vdd vdd in2 gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 vdd vdd clock_1/clkb vdd vdd vdd in3 gnd capacitors_1
Xcapacitors_1_4 input2 vdd vdd clock_1/clk vdd vdd vdd in2 gnd capacitors_1
Xcapacitors_1_5 input2 vdd vdd clock_1/clk vdd vdd vdd in3 gnd capacitors_1
Xcapacitors_1_6 input1 vdd vdd clock_1/clkb vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_7 input1 vdd vdd clock_1/clkb vdd vdd vdd in5 gnd capacitors_1
Xcapacitors_1_8 input1 vdd vdd clock_1/clkb vdd vdd vdd in6 gnd capacitors_1
Xcapacitors_1_9 input1 vdd vdd clock_1/clkb vdd vdd vdd in7 gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 vdd vdd clock_1/clk vdd vdd vdd in7 gnd capacitors_1
Xcapacitors_1_11 input2 vdd vdd clock_1/clk vdd vdd vdd in6 gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 vdd vdd clock_1/clk vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_12 input2 vdd vdd clock_1/clk vdd vdd vdd in5 gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clock_1/clk input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clock_1/clkb input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 m1_12464_n576# clock_1/clk 2.140857f
C1 input2 input1 3.059187f
C2 clock_1/clkb m1_12464_n576# 2.29778f
C3 vdd clock_1/clk 28.684513f
C4 vdd clock_1/clkb 32.261925f
C5 vdd input1 26.538095f
C6 vdd nmos_dnw3_0/vs 9.238383f
C7 clock_1/clkb nmos_dnw3_0/vs 2.218511f
C8 vdd input2 26.54464f
C9 input1 gnd 31.198782f
C10 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.396567f
C11 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079662f
C12 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634299f
C13 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398093f
C14 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.080289f
C15 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633591f
C16 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.392522f
C17 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079402f
C18 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634253f
C19 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398324f
C20 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079739f
C21 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633955f
C22 m1_4341_n519# gnd 3.765437f
C23 input2 gnd 30.578617f
C24 m1_12659_300# gnd 3.025714f
C25 m1_12464_n576# gnd 5.503336f
C26 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.397358f
C27 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079556f
C28 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634405f
C29 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.394424f
C30 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079656f
C31 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634067f
C32 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393486f
C33 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079731f
C34 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633915f
C35 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39339f
C36 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.07982f
C37 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633871f
C38 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.398049f
C39 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079472f
C40 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633938f
C41 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.396035f
C42 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079795f
C43 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634021f
C44 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.395022f
C45 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079731f
C46 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.634052f
C47 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.392135f
C48 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.078753f
C49 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.633513f
C50 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.338151f
C51 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.97841f
C52 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61055f
C53 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.33782f
C54 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.978384f
C55 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.610197f
C56 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.393725f
C57 clock_1/clk gnd 96.75779f
C58 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.080708f
C59 capacitor_8_1/capacitor_7_0/buffer_digital_0/in gnd 2.639487f
C60 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.397516f
C61 clock_1/clkb gnd 0.104535p
C62 vdd gnd 0.659544p
C63 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.079217f
C64 capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.639594f
C65 clock_1/a_2432_n962# gnd 8.693805f **FLOATING
C66 clock_1/a_2020_n482# gnd 2.56615f **FLOATING
C67 clock_1/a_344_102# gnd 2.809951f
C68 clock_1/a_2402_572# gnd 2.172722f
C69 clock_1/a_344_n986# gnd 2.381627f
C70 clock_1/a_3246_118# gnd 6.834443f
C71 nmos_dnw3_0/vs gnd 10.39343f
.ends

.subckt CP1_5_stage charge_pump1_2/in6 charge_pump1_2/in1 charge_pump1_2/in5 charge_pump1_2/vdd
+ charge_pump1_2/in4 charge_pump1_0/vin charge_pump1_2/in8 charge_pump1_2/m1_12464_n576#
+ charge_pump1_2/in3 charge_pump1_reverse_0/nmos_dnw3_0/vs charge_pump1_1/vin charge_pump1_2/gnd
+ buffer_digital_0/i charge_pump1_2/in2 charge_pump1_2/in7 charge_pump1_reverse_1/nmos_dnw3_0/vs
+ charge_pump1_2/vin
Xcharge_pump1_0 buffer_digital_0/i charge_pump1_0/input1 charge_pump1_0/input2 charge_pump1_2/vdd
+ charge_pump1_2/in1 charge_pump1_2/in2 charge_pump1_2/in6 charge_pump1_2/in7 charge_pump1_0/g1
+ charge_pump1_0/g2 charge_pump1_0/clk charge_pump1_0/clkb charge_pump1_reverse_0/nmos_dnw3_0/vs
+ charge_pump1_2/gnd charge_pump1_2/in4 charge_pump1_2/gnd charge_pump1_2/in3 charge_pump1_2/in5
+ charge_pump1_2/in8 charge_pump1_0/vin charge_pump1
Xcharge_pump1_1 charge_pump1_1/clk_in charge_pump1_1/input1 charge_pump1_1/input2
+ charge_pump1_2/vdd charge_pump1_2/in1 charge_pump1_2/in2 charge_pump1_2/in6 charge_pump1_2/in7
+ charge_pump1_1/g1 charge_pump1_1/g2 charge_pump1_1/clk charge_pump1_1/clkb charge_pump1_reverse_1/nmos_dnw3_0/vs
+ charge_pump1_1/a_3340_18086# charge_pump1_2/in4 charge_pump1_2/gnd charge_pump1_2/in3
+ charge_pump1_2/in5 charge_pump1_2/in8 charge_pump1_1/vin charge_pump1
Xcharge_pump1_2 charge_pump1_2/clk_in charge_pump1_2/input1 charge_pump1_2/input2
+ charge_pump1_2/vdd charge_pump1_2/in1 charge_pump1_2/in2 charge_pump1_2/in6 charge_pump1_2/in7
+ charge_pump1_2/g1 charge_pump1_2/g2 charge_pump1_2/clk charge_pump1_2/clkb charge_pump1_2/m1_12464_n576#
+ charge_pump1_2/a_3340_18086# charge_pump1_2/in4 charge_pump1_2/gnd charge_pump1_2/in3
+ charge_pump1_2/in5 charge_pump1_2/in8 charge_pump1_2/vin charge_pump1
Xcharge_pump1_reverse_0 charge_pump1_reverse_0/input1 charge_pump1_reverse_0/input2
+ charge_pump1_2/in8 charge_pump1_2/in7 charge_pump1_2/in3 charge_pump1_2/in2 charge_pump1_2/vdd
+ charge_pump1_1/vin buffer_digital_1/in charge_pump1_2/gnd charge_pump1_2/gnd charge_pump1_2/in5
+ charge_pump1_2/in6 charge_pump1_2/in4 charge_pump1_2/in1 charge_pump1_reverse_0/nmos_dnw3_0/vs
+ charge_pump1_reverse
Xbuffer_digital_0 buffer_digital_0/i buffer_digital_1/i charge_pump1_2/vdd charge_pump1_2/gnd
+ buffer_digital_0/a_116_148# buffer_digital
Xcharge_pump1_reverse_1 charge_pump1_reverse_1/input1 charge_pump1_reverse_1/input2
+ charge_pump1_2/in8 charge_pump1_2/in7 charge_pump1_2/in3 charge_pump1_2/in2 charge_pump1_2/vdd
+ charge_pump1_2/vin charge_pump1_reverse_1/clock_1/clk_in charge_pump1_2/gnd charge_pump1_2/gnd
+ charge_pump1_2/in5 charge_pump1_2/in6 charge_pump1_2/in4 charge_pump1_2/in1 charge_pump1_reverse_1/nmos_dnw3_0/vs
+ charge_pump1_reverse
Xbuffer_digital_1 buffer_digital_1/i buffer_digital_1/in charge_pump1_2/vdd charge_pump1_2/gnd
+ m1_30262_n2398# buffer_digital
X0 a_73934_n2624# charge_pump1_1/clk_in charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X1 a_100152_n2424# a_99934_n2424# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X2 charge_pump1_reverse_1/clock_1/clk_in a_80522_n2634# charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X3 charge_pump1_reverse_1/clock_1/clk_in a_80522_n2634# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X4 a_48152_n2524# a_47934_n2524# charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X5 a_54522_n2534# a_48152_n2524# charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X6 a_48152_n2524# a_47934_n2524# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X7 a_54522_n2534# a_48152_n2524# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X8 a_106522_n2434# a_100152_n2424# charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X9 a_47934_n2524# buffer_digital_1/in charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X10 a_106522_n2434# a_100152_n2424# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X11 a_47934_n2524# buffer_digital_1/in charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X12 charge_pump1_1/clk_in a_54522_n2534# charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X13 charge_pump1_1/clk_in a_54522_n2534# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X14 a_74152_n2624# a_73934_n2624# charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X15 a_80522_n2634# a_74152_n2624# charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X16 charge_pump1_2/clk_in a_106522_n2434# charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X17 a_74152_n2624# a_73934_n2624# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X18 a_80522_n2634# a_74152_n2624# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X19 a_99934_n2424# charge_pump1_reverse_1/clock_1/clk_in charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X20 charge_pump1_2/clk_in a_106522_n2434# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X21 a_99934_n2424# charge_pump1_reverse_1/clock_1/clk_in charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.3654 pd=3.1 as=0.3654 ps=3.1 w=1.26 l=0.15
X22 a_100152_n2424# a_99934_n2424# charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X23 a_73934_n2624# charge_pump1_1/clk_in charge_pump1_2/gnd charge_pump1_2/gnd sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
C0 buffer_digital_0/i charge_pump1_2/vdd 4.615536f
C1 charge_pump1_2/vdd charge_pump1_2/in5 3.750112f
C2 charge_pump1_2/vdd charge_pump1_reverse_1/clock_1/clk_in 5.607365f
C3 charge_pump1_2/vdd buffer_digital_1/in 4.877749f
C4 charge_pump1_2/vdd charge_pump1_2/in3 3.749226f
C5 charge_pump1_2/vdd charge_pump1_2/in7 3.658818f
C6 charge_pump1_2/vdd charge_pump1_1/clk_in 5.599668f
C7 charge_pump1_2/vdd charge_pump1_2/in1 3.688278f
C8 charge_pump1_2/vdd charge_pump1_2/in2 3.748251f
C9 charge_pump1_2/vdd charge_pump1_2/in6 3.780672f
C10 charge_pump1_2/vdd charge_pump1_2/in8 3.690953f
C11 charge_pump1_2/vdd charge_pump1_2/clk_in 2.833448f
C12 charge_pump1_2/vdd charge_pump1_2/in4 3.75142f
C13 a_100152_n2424# charge_pump1_2/gnd 2.75745f
C14 a_74152_n2624# charge_pump1_2/gnd 2.81589f
C15 a_48152_n2524# charge_pump1_2/gnd 2.95405f
C16 charge_pump1_reverse_1/input1 charge_pump1_2/gnd 22.596436f
C17 charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C18 charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C19 charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C20 charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C21 charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C22 charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C23 charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C24 charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C25 charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C26 charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C27 charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C28 charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C29 charge_pump1_reverse_1/m1_4341_n519# charge_pump1_2/gnd 3.33176f
C30 charge_pump1_reverse_1/input2 charge_pump1_2/gnd 22.21436f
C31 charge_pump1_reverse_1/m1_12659_300# charge_pump1_2/gnd 2.683598f
C32 charge_pump1_2/vin charge_pump1_2/gnd 14.30258f
C33 charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C34 charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C35 charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C36 charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C37 charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C38 charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C39 charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C40 charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C41 charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C42 charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C43 charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C44 charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C45 charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C46 charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C47 charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C48 charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C49 charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C50 charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C51 charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C52 charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C53 charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C54 charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C55 charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C56 charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C57 charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C58 charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C59 charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C60 charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C61 charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C62 charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C63 charge_pump1_2/in8 charge_pump1_2/gnd 10.682923f
C64 charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C65 charge_pump1_reverse_1/clock_1/clk charge_pump1_2/gnd 94.62247f
C66 charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C67 charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C68 charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C69 charge_pump1_reverse_1/clock_1/clkb charge_pump1_2/gnd 0.1013p
C70 charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C71 charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C72 charge_pump1_reverse_1/clock_1/a_2432_n962# charge_pump1_2/gnd 8.68424f **FLOATING
C73 charge_pump1_reverse_1/clock_1/a_2020_n482# charge_pump1_2/gnd 2.56615f **FLOATING
C74 charge_pump1_reverse_1/clock_1/a_344_102# charge_pump1_2/gnd 2.809951f
C75 charge_pump1_reverse_1/clock_1/a_2402_572# charge_pump1_2/gnd 2.172722f
C76 charge_pump1_reverse_1/clock_1/a_344_n986# charge_pump1_2/gnd 2.381627f
C77 charge_pump1_reverse_1/clock_1/clk_in charge_pump1_2/gnd 16.46123f
C78 charge_pump1_reverse_1/clock_1/a_3246_118# charge_pump1_2/gnd 6.834443f
C79 buffer_digital_1/i charge_pump1_2/gnd 2.551267f
C80 charge_pump1_reverse_0/input1 charge_pump1_2/gnd 22.596436f
C81 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C82 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C83 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C84 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C85 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C86 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C87 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C88 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C89 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C90 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C91 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C92 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C93 charge_pump1_reverse_0/m1_4341_n519# charge_pump1_2/gnd 3.33176f
C94 charge_pump1_reverse_0/input2 charge_pump1_2/gnd 22.21436f
C95 charge_pump1_reverse_0/m1_12659_300# charge_pump1_2/gnd 2.683598f
C96 charge_pump1_1/vin charge_pump1_2/gnd 14.23653f
C97 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C98 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C99 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C100 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C101 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C102 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C103 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C104 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C105 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C106 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C107 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C108 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C109 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C110 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C111 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C112 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C113 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C114 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C115 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C116 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C117 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C118 charge_pump1_2/in6 charge_pump1_2/gnd 10.482664f
C119 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C120 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C121 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C122 charge_pump1_2/in7 charge_pump1_2/gnd 10.354812f
C123 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C124 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C125 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C126 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C127 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C128 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C129 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C130 charge_pump1_reverse_0/clock_1/clk charge_pump1_2/gnd 94.59402f
C131 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C132 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C133 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C134 charge_pump1_reverse_0/clock_1/clkb charge_pump1_2/gnd 0.101491p
C135 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C136 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C137 charge_pump1_reverse_0/clock_1/a_2432_n962# charge_pump1_2/gnd 8.68424f **FLOATING
C138 charge_pump1_reverse_0/clock_1/a_2020_n482# charge_pump1_2/gnd 2.56615f **FLOATING
C139 charge_pump1_reverse_0/clock_1/a_344_102# charge_pump1_2/gnd 2.809951f
C140 charge_pump1_reverse_0/clock_1/a_2402_572# charge_pump1_2/gnd 2.172722f
C141 charge_pump1_reverse_0/clock_1/a_344_n986# charge_pump1_2/gnd 2.381627f
C142 buffer_digital_1/in charge_pump1_2/gnd 13.948167f
C143 charge_pump1_reverse_0/clock_1/a_3246_118# charge_pump1_2/gnd 6.834443f
C144 charge_pump1_2/a_3340_18086# charge_pump1_2/gnd 6.04146f
C145 charge_pump1_2/input1 charge_pump1_2/gnd 22.463037f
C146 charge_pump1_2/input2 charge_pump1_2/gnd 22.175129f
C147 charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C148 charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C149 charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C150 charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C151 charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C152 charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C153 charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C154 charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C155 charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C156 charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C157 charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C158 charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C159 charge_pump1_2/m1_4341_n519# charge_pump1_2/gnd 3.771611f
C160 charge_pump1_2/m1_12659_300# charge_pump1_2/gnd 2.538747f
C161 charge_pump1_2/m1_12464_n576# charge_pump1_2/gnd 4.258816f
C162 charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C163 charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C164 charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C165 charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C166 charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C167 charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C168 charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C169 charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C170 charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C171 charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C172 charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C173 charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C174 charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C175 charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C176 charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C177 charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C178 charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C179 charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C180 charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C181 charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C182 charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C183 charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C184 charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C185 charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C186 charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C187 charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C188 charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C189 charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C190 charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C191 charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C192 charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C193 charge_pump1_2/clkb charge_pump1_2/gnd 89.87499f
C194 charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C195 charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C196 charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C197 charge_pump1_2/clk charge_pump1_2/gnd 89.19299f
C198 charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C199 charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C200 charge_pump1_2/clock_0/a_2432_n962# charge_pump1_2/gnd 8.68424f **FLOATING
C201 charge_pump1_2/clock_0/a_2020_n482# charge_pump1_2/gnd 2.56615f **FLOATING
C202 charge_pump1_2/clock_0/a_344_102# charge_pump1_2/gnd 2.809951f
C203 charge_pump1_2/clock_0/a_2402_572# charge_pump1_2/gnd 2.172722f
C204 charge_pump1_2/clock_0/a_344_n986# charge_pump1_2/gnd 2.381627f
C205 charge_pump1_2/clk_in charge_pump1_2/gnd 11.703724f
C206 charge_pump1_2/clock_0/a_3246_118# charge_pump1_2/gnd 6.834443f
C207 charge_pump1_2/g2 charge_pump1_2/gnd 2.344427f
C208 charge_pump1_1/a_3340_18086# charge_pump1_2/gnd 6.141427f
C209 charge_pump1_1/input1 charge_pump1_2/gnd 22.463037f
C210 charge_pump1_1/input2 charge_pump1_2/gnd 22.175129f
C211 charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C212 charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C213 charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C214 charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C215 charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C216 charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C217 charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C218 charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C219 charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C220 charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C221 charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C222 charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C223 charge_pump1_1/m1_4341_n519# charge_pump1_2/gnd 3.771611f
C224 charge_pump1_1/m1_12659_300# charge_pump1_2/gnd 2.538747f
C225 charge_pump1_reverse_1/nmos_dnw3_0/vs charge_pump1_2/gnd 14.559652f
C226 charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C227 charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C228 charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C229 charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C230 charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C231 charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C232 charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C233 charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C234 charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C235 charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C236 charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C237 charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C238 charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C239 charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C240 charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C241 charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C242 charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C243 charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C244 charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C245 charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C246 charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C247 charge_pump1_2/in3 charge_pump1_2/gnd 10.433572f
C248 charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C249 charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C250 charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C251 charge_pump1_2/in2 charge_pump1_2/gnd 10.455082f
C252 charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C253 charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C254 charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C255 charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C256 charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C257 charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C258 charge_pump1_2/in1 charge_pump1_2/gnd 9.979585f
C259 charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C260 charge_pump1_1/clkb charge_pump1_2/gnd 89.84497f
C261 charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C262 charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C263 charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C264 charge_pump1_1/clk charge_pump1_2/gnd 89.19739f
C265 charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C266 charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C267 charge_pump1_1/clock_0/a_2432_n962# charge_pump1_2/gnd 8.68424f **FLOATING
C268 charge_pump1_1/clock_0/a_2020_n482# charge_pump1_2/gnd 2.56615f **FLOATING
C269 charge_pump1_1/clock_0/a_344_102# charge_pump1_2/gnd 2.809951f
C270 charge_pump1_1/clock_0/a_2402_572# charge_pump1_2/gnd 2.172722f
C271 charge_pump1_1/clock_0/a_344_n986# charge_pump1_2/gnd 2.381627f
C272 charge_pump1_1/clk_in charge_pump1_2/gnd 19.857828f
C273 charge_pump1_1/clock_0/a_3246_118# charge_pump1_2/gnd 6.834443f
C274 charge_pump1_1/g2 charge_pump1_2/gnd 2.344427f
C275 charge_pump1_0/input1 charge_pump1_2/gnd 22.463037f
C276 charge_pump1_0/input2 charge_pump1_2/gnd 22.175129f
C277 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C278 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C279 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C280 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C281 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C282 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C283 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C284 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C285 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C286 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C287 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C288 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C289 charge_pump1_0/m1_4341_n519# charge_pump1_2/gnd 3.771611f
C290 charge_pump1_0/m1_12659_300# charge_pump1_2/gnd 2.538747f
C291 charge_pump1_reverse_0/nmos_dnw3_0/vs charge_pump1_2/gnd 14.770787f
C292 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C293 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C294 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C295 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C296 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C297 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C298 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C299 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C300 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C301 charge_pump1_2/in5 charge_pump1_2/gnd 10.548278f
C302 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C303 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C304 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C305 charge_pump1_2/in4 charge_pump1_2/gnd 10.550569f
C306 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C307 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C308 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C309 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C310 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C311 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C312 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C313 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C314 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C315 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C316 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C317 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C318 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C319 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C320 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C321 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C322 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C323 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C324 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C325 charge_pump1_0/clkb charge_pump1_2/gnd 89.96071f
C326 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C327 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C328 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump1_2/gnd 2.337696f
C329 charge_pump1_0/clk charge_pump1_2/gnd 89.28753f
C330 charge_pump1_2/vdd charge_pump1_2/gnd 2.526324p
C331 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump1_2/gnd 9.978376f
C332 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in charge_pump1_2/gnd 2.608221f
C333 charge_pump1_0/clock_0/a_2432_n962# charge_pump1_2/gnd 8.68424f **FLOATING
C334 charge_pump1_0/clock_0/a_2020_n482# charge_pump1_2/gnd 2.56615f **FLOATING
C335 charge_pump1_0/clock_0/a_344_102# charge_pump1_2/gnd 2.809951f
C336 charge_pump1_0/clock_0/a_2402_572# charge_pump1_2/gnd 2.172722f
C337 charge_pump1_0/clock_0/a_344_n986# charge_pump1_2/gnd 2.381627f
C338 buffer_digital_0/i charge_pump1_2/gnd 23.756302f
C339 charge_pump1_0/clock_0/a_3246_118# charge_pump1_2/gnd 6.834443f
C340 charge_pump1_0/g2 charge_pump1_2/gnd 2.344427f
C341 charge_pump1_0/vin charge_pump1_2/gnd 10.369197f
.ends

.subckt reconfigurable_CP_lvs1
XCP2_5_stage_1 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/vs CP2_5_stage_1/buffer_digital_7/in
+ CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/out2 CP2_5_stage_1/charge_pump_2/out
+ CP2_5_stage_1/charge_pump_0/out CP1_5_stage_0/charge_pump1_2/vdd CP2_5_stage_1/charge_pump_2/in3
+ CP2_5_stage_1/charge_pump_0/vin CP2_5_stage_1/charge_pump_2/in4 CP2_5_stage_1/charge_pump_reverse_1/clock_0/clk
+ CP2_5_stage_1/charge_pump_0/vs CP2_5_stage_1/buffer_digital_4/i CP2_5_stage_1/charge_pump_2/in5
+ CP2_5_stage_1/charge_pump_2/in6 CP2_5_stage_1/charge_pump_1/vs CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/vs
+ CP2_5_stage_1/charge_pump_2/in8 CP2_5_stage_1/charge_pump_2/in1 CP2_5_stage_1/buffer_digital_0/i
+ CP2_5_stage_1/buffer_digital_6/i VSUBS CP2_5_stage_1/charge_pump_2/in7 CP2_5_stage_1/charge_pump_2/vs
+ CP2_5_stage_1/charge_pump_2/in2 CP2_5_stage
XCP2_5_stage_0 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/vs CP2_5_stage_1/buffer_digital_0/i
+ VSUBS CP2_5_stage_1/charge_pump_0/vin CP2_5_stage_0/charge_pump_0/out CP1_5_stage_0/charge_pump1_2/vdd
+ CP2_5_stage_1/charge_pump_2/in6 CP2_5_stage_0/charge_pump_0/vin CP2_5_stage_1/charge_pump_2/in5
+ VSUBS CP2_5_stage_0/charge_pump_0/vs CP2_5_stage_0/buffer_digital_4/i CP2_5_stage_1/charge_pump_2/in4
+ CP2_5_stage_1/charge_pump_2/in3 CP2_5_stage_0/charge_pump_1/vs CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/vs
+ CP2_5_stage_1/charge_pump_2/in1 CP2_5_stage_1/charge_pump_2/in8 CP2_5_stage_0/buffer_digital_0/i
+ CP2_5_stage_0/buffer_digital_6/i VSUBS CP2_5_stage_1/charge_pump_2/in2 CP2_5_stage_0/charge_pump_2/vs
+ CP2_5_stage_1/charge_pump_2/in7 CP2_5_stage
XCP1_5_stage_0 CP2_5_stage_1/charge_pump_2/in6 CP2_5_stage_1/charge_pump_2/in1 CP2_5_stage_1/charge_pump_2/in5
+ CP1_5_stage_0/charge_pump1_2/vdd CP2_5_stage_1/charge_pump_2/in4 CP1_5_stage_0/charge_pump1_0/vin
+ CP2_5_stage_1/charge_pump_2/in8 m2_128295_42196# CP2_5_stage_1/charge_pump_2/in3
+ CP1_5_stage_0/charge_pump1_reverse_0/nmos_dnw3_0/vs CP1_5_stage_0/charge_pump1_1/vin
+ VSUBS CP2_5_stage_1/buffer_digital_0/i CP2_5_stage_1/charge_pump_2/in2 CP2_5_stage_1/charge_pump_2/in7
+ CP1_5_stage_0/charge_pump1_reverse_1/nmos_dnw3_0/vs CP1_5_stage_0/charge_pump1_2/vin
+ CP1_5_stage
C0 CP2_5_stage_1/charge_pump_2/in1 CP2_5_stage_1/charge_pump_2/in8 3.24343f
C1 CP2_5_stage_1/charge_pump_2/in6 CP2_5_stage_1/charge_pump_2/in5 9.099842f
C2 CP2_5_stage_1/charge_pump_2/in7 CP2_5_stage_1/charge_pump_2/in8 5.41224f
C3 CP2_5_stage_1/charge_pump_2/in4 CP2_5_stage_1/charge_pump_2/in5 10.4178f
C4 CP2_5_stage_1/charge_pump_2/in3 CP2_5_stage_1/charge_pump_2/in4 9.06413f
C5 CP2_5_stage_1/charge_pump_2/in7 CP2_5_stage_1/charge_pump_2/in6 8.147181f
C6 CP2_5_stage_1/charge_pump_2/in2 CP2_5_stage_1/buffer_digital_0/i 2.278516f
C7 CP2_5_stage_1/charge_pump_2/in7 CP2_5_stage_1/charge_pump_2/in3 2.23645f
C8 CP2_5_stage_1/charge_pump_2/in2 CP2_5_stage_1/charge_pump_2/in3 8.175771f
C9 CP2_5_stage_1/charge_pump_2/in1 CP2_5_stage_1/charge_pump_2/in2 13.3543f
C10 CP2_5_stage_1/charge_pump_2/in7 CP2_5_stage_1/charge_pump_2/in2 2.68839f
C11 CP1_5_stage_0/charge_pump1_2/vdd CP2_5_stage_1/buffer_digital_0/i 2.997349f
C12 CP1_5_stage_0/a_100152_n2424# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.75745f **FLOATING
C13 CP1_5_stage_0/a_74152_n2624# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.81589f **FLOATING
C14 CP1_5_stage_0/a_48152_n2524# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.95405f **FLOATING
C15 CP1_5_stage_0/charge_pump1_reverse_1/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.596436f
C16 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C17 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C18 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C19 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C20 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C21 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C22 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C23 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C24 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C25 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C26 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C27 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C28 CP1_5_stage_0/charge_pump1_reverse_1/m1_4341_n519# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 3.33176f
C29 CP1_5_stage_0/charge_pump1_reverse_1/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.21436f
C30 CP1_5_stage_0/charge_pump1_reverse_1/m1_12659_300# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.683598f
C31 CP1_5_stage_0/charge_pump1_2/vin CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.262471f
C32 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C33 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C34 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C35 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C36 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C37 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C38 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C39 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C40 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C41 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C42 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C43 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C44 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C45 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C46 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C47 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C48 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C49 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C50 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C51 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C52 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C53 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C54 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C55 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C56 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C57 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C58 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C59 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C60 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C61 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C62 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C63 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 94.613235f
C64 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C65 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C66 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C67 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 0.10133p
C68 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C69 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C70 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C71 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C72 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C73 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C74 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C75 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/clk_in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 16.172987f
C76 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C77 CP1_5_stage_0/buffer_digital_1/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.523045f
C78 CP1_5_stage_0/charge_pump1_reverse_0/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.596436f
C79 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C80 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C81 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C82 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C83 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C84 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C85 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C86 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C87 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C88 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C89 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C90 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C91 CP1_5_stage_0/charge_pump1_reverse_0/m1_4341_n519# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 3.33176f
C92 CP1_5_stage_0/charge_pump1_reverse_0/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.21436f
C93 CP1_5_stage_0/charge_pump1_reverse_0/m1_12659_300# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.683598f
C94 CP1_5_stage_0/charge_pump1_1/vin CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.201631f
C95 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C96 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C97 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C98 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C99 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C100 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C101 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C102 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C103 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C104 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C105 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C106 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C107 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C108 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C109 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C110 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C111 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C112 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C113 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C114 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C115 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C116 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C117 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C118 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C119 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C120 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C121 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C122 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C123 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C124 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C125 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C126 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 94.613235f
C127 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C128 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C129 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C130 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 0.10133p
C131 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C132 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C133 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C134 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C135 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C136 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C137 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C138 CP1_5_stage_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 13.623026f
C139 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C140 CP1_5_stage_0/charge_pump1_2/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.463037f
C141 CP1_5_stage_0/charge_pump1_2/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.175129f
C142 CP1_5_stage_0/charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C143 CP1_5_stage_0/charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C144 CP1_5_stage_0/charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C145 CP1_5_stage_0/charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C146 CP1_5_stage_0/charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C147 CP1_5_stage_0/charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C148 CP1_5_stage_0/charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C149 CP1_5_stage_0/charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C150 CP1_5_stage_0/charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C151 CP1_5_stage_0/charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C152 CP1_5_stage_0/charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C153 CP1_5_stage_0/charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C154 CP1_5_stage_0/charge_pump1_2/m1_4341_n519# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 3.771611f
C155 CP1_5_stage_0/charge_pump1_2/m1_12659_300# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.538747f
C156 m2_128295_42196# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.524068f
C157 CP1_5_stage_0/charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C158 CP1_5_stage_0/charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C159 CP1_5_stage_0/charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C160 CP1_5_stage_0/charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C161 CP1_5_stage_0/charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C162 CP1_5_stage_0/charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C163 CP1_5_stage_0/charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C164 CP1_5_stage_0/charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C165 CP1_5_stage_0/charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C166 CP1_5_stage_0/charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C167 CP1_5_stage_0/charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C168 CP1_5_stage_0/charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C169 CP1_5_stage_0/charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C170 CP1_5_stage_0/charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C171 CP1_5_stage_0/charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C172 CP1_5_stage_0/charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C173 CP1_5_stage_0/charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C174 CP1_5_stage_0/charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C175 CP1_5_stage_0/charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C176 CP1_5_stage_0/charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C177 CP1_5_stage_0/charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C178 CP1_5_stage_0/charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C179 CP1_5_stage_0/charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C180 CP1_5_stage_0/charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C181 CP1_5_stage_0/charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C182 CP1_5_stage_0/charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C183 CP1_5_stage_0/charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C184 CP1_5_stage_0/charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C185 CP1_5_stage_0/charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C186 CP1_5_stage_0/charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C187 CP1_5_stage_0/charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C188 CP1_5_stage_0/charge_pump1_2/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 89.87449f
C189 CP1_5_stage_0/charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C190 CP1_5_stage_0/charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C191 CP1_5_stage_0/charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C192 CP1_5_stage_0/charge_pump1_2/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 89.042244f
C193 CP1_5_stage_0/charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C194 CP1_5_stage_0/charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C195 CP1_5_stage_0/charge_pump1_2/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C196 CP1_5_stage_0/charge_pump1_2/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C197 CP1_5_stage_0/charge_pump1_2/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C198 CP1_5_stage_0/charge_pump1_2/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C199 CP1_5_stage_0/charge_pump1_2/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C200 CP1_5_stage_0/charge_pump1_2/clk_in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 11.702157f
C201 CP1_5_stage_0/charge_pump1_2/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C202 CP1_5_stage_0/charge_pump1_2/g2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.344427f
C203 CP1_5_stage_0/charge_pump1_1/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.463037f
C204 CP1_5_stage_0/charge_pump1_1/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.175129f
C205 CP1_5_stage_0/charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C206 CP1_5_stage_0/charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C207 CP1_5_stage_0/charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C208 CP1_5_stage_0/charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C209 CP1_5_stage_0/charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C210 CP1_5_stage_0/charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C211 CP1_5_stage_0/charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C212 CP1_5_stage_0/charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C213 CP1_5_stage_0/charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C214 CP1_5_stage_0/charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C215 CP1_5_stage_0/charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C216 CP1_5_stage_0/charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C217 CP1_5_stage_0/charge_pump1_1/m1_4341_n519# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 3.771611f
C218 CP1_5_stage_0/charge_pump1_1/m1_12659_300# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.538747f
C219 CP1_5_stage_0/charge_pump1_reverse_1/nmos_dnw3_0/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.50642f
C220 CP1_5_stage_0/charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C221 CP1_5_stage_0/charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C222 CP1_5_stage_0/charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C223 CP1_5_stage_0/charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C224 CP1_5_stage_0/charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C225 CP1_5_stage_0/charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C226 CP1_5_stage_0/charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C227 CP1_5_stage_0/charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C228 CP1_5_stage_0/charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C229 CP1_5_stage_0/charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C230 CP1_5_stage_0/charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C231 CP1_5_stage_0/charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C232 CP1_5_stage_0/charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C233 CP1_5_stage_0/charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C234 CP1_5_stage_0/charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C235 CP1_5_stage_0/charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C236 CP1_5_stage_0/charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C237 CP1_5_stage_0/charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C238 CP1_5_stage_0/charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C239 CP1_5_stage_0/charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C240 CP1_5_stage_0/charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C241 CP1_5_stage_0/charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C242 CP1_5_stage_0/charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C243 CP1_5_stage_0/charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C244 CP1_5_stage_0/charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C245 CP1_5_stage_0/charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C246 CP1_5_stage_0/charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C247 CP1_5_stage_0/charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C248 CP1_5_stage_0/charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C249 CP1_5_stage_0/charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C250 CP1_5_stage_0/charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C251 CP1_5_stage_0/charge_pump1_1/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 89.87499f
C252 CP1_5_stage_0/charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C253 CP1_5_stage_0/charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C254 CP1_5_stage_0/charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C255 CP1_5_stage_0/charge_pump1_1/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 89.042244f
C256 CP1_5_stage_0/charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C257 CP1_5_stage_0/charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C258 CP1_5_stage_0/charge_pump1_1/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C259 CP1_5_stage_0/charge_pump1_1/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C260 CP1_5_stage_0/charge_pump1_1/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C261 CP1_5_stage_0/charge_pump1_1/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C262 CP1_5_stage_0/charge_pump1_1/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C263 CP1_5_stage_0/charge_pump1_1/clk_in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 19.85626f
C264 CP1_5_stage_0/charge_pump1_1/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C265 CP1_5_stage_0/charge_pump1_1/g2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.344427f
C266 CP1_5_stage_0/charge_pump1_0/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.463037f
C267 CP1_5_stage_0/charge_pump1_0/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 22.175129f
C268 CP1_5_stage_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C269 CP1_5_stage_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C270 CP1_5_stage_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C271 CP1_5_stage_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C272 CP1_5_stage_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C273 CP1_5_stage_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C274 CP1_5_stage_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C275 CP1_5_stage_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C276 CP1_5_stage_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C277 CP1_5_stage_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C278 CP1_5_stage_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C279 CP1_5_stage_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C280 CP1_5_stage_0/charge_pump1_0/m1_4341_n519# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 3.771611f
C281 CP1_5_stage_0/charge_pump1_0/m1_12659_300# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.538747f
C282 CP1_5_stage_0/charge_pump1_reverse_0/nmos_dnw3_0/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.690079f
C283 CP1_5_stage_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C284 CP1_5_stage_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C285 CP1_5_stage_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C286 CP1_5_stage_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C287 CP1_5_stage_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C288 CP1_5_stage_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C289 CP1_5_stage_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C290 CP1_5_stage_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C291 CP1_5_stage_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C292 CP1_5_stage_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C293 CP1_5_stage_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C294 CP1_5_stage_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C295 CP1_5_stage_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C296 CP1_5_stage_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C297 CP1_5_stage_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C298 CP1_5_stage_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C299 CP1_5_stage_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C300 CP1_5_stage_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C301 CP1_5_stage_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C302 CP1_5_stage_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C303 CP1_5_stage_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608206f
C304 CP1_5_stage_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C305 CP1_5_stage_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C306 CP1_5_stage_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C307 CP1_5_stage_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C308 CP1_5_stage_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C309 CP1_5_stage_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C310 CP1_5_stage_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C311 CP1_5_stage_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C312 CP1_5_stage_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C313 CP1_5_stage_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C314 CP1_5_stage_0/charge_pump1_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 89.87499f
C315 CP1_5_stage_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C316 CP1_5_stage_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C317 CP1_5_stage_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C318 CP1_5_stage_0/charge_pump1_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 89.017944f
C319 CP1_5_stage_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C320 CP1_5_stage_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.608221f
C321 CP1_5_stage_0/charge_pump1_0/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C322 CP1_5_stage_0/charge_pump1_0/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C323 CP1_5_stage_0/charge_pump1_0/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C324 CP1_5_stage_0/charge_pump1_0/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C325 CP1_5_stage_0/charge_pump1_0/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C326 CP1_5_stage_0/charge_pump1_0/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C327 CP1_5_stage_0/charge_pump1_0/g2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.344427f
C328 CP1_5_stage_0/charge_pump1_0/vin CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 10.366855f
C329 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.79532f
C330 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C331 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C332 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C333 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C334 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C335 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C336 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.234749f
C337 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C338 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C339 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C340 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C341 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C342 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C343 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C344 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C345 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C346 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C347 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C348 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C349 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C350 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C351 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C352 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/out1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.749125f
C353 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C354 CP2_5_stage_0/charge_pump_reverse_1/clock_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 91.59107f
C355 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C356 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C357 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C358 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C359 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C360 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C361 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C362 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C363 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C364 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C365 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C366 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C367 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C368 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C369 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C370 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C371 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C372 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C373 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C374 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C375 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C376 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C377 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C378 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C379 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C380 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C381 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C382 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C383 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C384 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C385 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C386 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C387 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.425359f
C388 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.79532f
C389 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C390 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C391 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C392 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C393 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C394 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C395 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.234749f
C396 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C397 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C398 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C399 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C400 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C401 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C402 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C403 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C404 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C405 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C406 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C407 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C408 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C409 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C410 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C411 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/out1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.791632f
C412 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C413 CP2_5_stage_0/charge_pump_reverse_0/clock_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 91.6145f
C414 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C415 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C416 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C417 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C418 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C419 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C420 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C421 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C422 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C423 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C424 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C425 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C426 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C427 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C428 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C429 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C430 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C431 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C432 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C433 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C434 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C435 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C436 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C437 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/out2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.939422f
C438 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C439 CP2_5_stage_0/charge_pump_reverse_0/clock_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 85.213036f
C440 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C441 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C442 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C443 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C444 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C445 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C446 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C447 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C448 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.425359f
C449 CP2_5_stage_0/buffer_digital_6/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 10.265736f
C450 CP2_5_stage_0/buffer_digital_2/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.585812f
C451 CP2_5_stage_0/charge_pump_2/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.962303f
C452 CP2_5_stage_0/charge_pump_2/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C453 CP2_5_stage_0/charge_pump_2/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C454 CP2_5_stage_0/charge_pump_2/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C455 CP2_5_stage_0/charge_pump_2/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C456 CP2_5_stage_0/charge_pump_2/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C457 CP2_5_stage_0/charge_pump_2/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C458 CP2_5_stage_0/charge_pump_2/g2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.457181f
C459 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C460 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C461 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C462 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C463 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C464 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C465 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C466 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C467 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C468 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C469 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C470 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C471 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C472 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C473 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C474 CP2_5_stage_0/charge_pump_2/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.031953f
C475 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C476 CP2_5_stage_0/charge_pump_2/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 82.335495f
C477 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C478 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C479 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C480 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C481 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C482 CP2_5_stage_1/charge_pump_2/in2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 32.59423f
C483 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C484 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C485 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C486 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C487 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C488 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C489 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C490 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C491 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C492 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C493 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C494 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C495 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C496 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C497 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C498 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C499 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C500 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C501 CP2_5_stage_0/charge_pump_2/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.390842f
C502 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C503 CP2_5_stage_0/charge_pump_2/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 83.99082f
C504 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C505 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C506 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C507 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C508 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C509 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C510 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C511 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C512 CP2_5_stage_0/charge_pump_2/g1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.656219f
C513 CP2_5_stage_0/buffer_digital_1/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.342446f
C514 CP2_5_stage_0/charge_pump_1/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.96237f
C515 CP2_5_stage_0/charge_pump_1/out CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 3.305988f
C516 CP2_5_stage_0/charge_pump_1/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C517 CP2_5_stage_0/charge_pump_1/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C518 CP2_5_stage_0/charge_pump_1/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C519 CP2_5_stage_0/charge_pump_1/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C520 CP2_5_stage_0/charge_pump_1/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C521 CP2_5_stage_0/buffer_digital_4/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.591777f
C522 CP2_5_stage_0/charge_pump_1/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C523 CP2_5_stage_0/charge_pump_1/g2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.514679f
C524 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C525 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C526 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C527 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C528 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C529 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C530 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C531 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C532 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C533 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C534 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C535 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C536 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C537 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C538 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C539 CP2_5_stage_0/charge_pump_1/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.031953f
C540 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C541 CP2_5_stage_0/charge_pump_1/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 82.33631f
C542 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C543 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C544 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C545 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C546 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C547 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C548 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C549 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C550 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C551 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C552 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C553 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C554 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C555 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C556 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C557 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C558 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C559 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C560 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C561 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C562 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C563 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C564 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C565 CP2_5_stage_0/charge_pump_1/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.390842f
C566 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C567 CP2_5_stage_0/charge_pump_1/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 84.10069f
C568 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C569 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C570 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C571 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C572 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C573 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C574 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C575 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C576 CP2_5_stage_0/charge_pump_1/g1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.656795f
C577 CP2_5_stage_0/charge_pump_0/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.96237f
C578 CP2_5_stage_0/charge_pump_0/out CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.12709f
C579 CP2_5_stage_0/charge_pump_0/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C580 CP2_5_stage_0/charge_pump_0/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C581 CP2_5_stage_0/charge_pump_0/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C582 CP2_5_stage_0/charge_pump_0/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C583 CP2_5_stage_0/charge_pump_0/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C584 CP2_5_stage_0/buffer_digital_0/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 17.01914f
C585 CP2_5_stage_0/charge_pump_0/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C586 CP2_5_stage_0/charge_pump_0/g2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.457593f
C587 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C588 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C589 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C590 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C591 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C592 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C593 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C594 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C595 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C596 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C597 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C598 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C599 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C600 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C601 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C602 CP2_5_stage_0/charge_pump_0/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.031953f
C603 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C604 CP2_5_stage_0/charge_pump_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 82.35288f
C605 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C606 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C607 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C608 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C609 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C610 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C611 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C612 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C613 CP2_5_stage_1/charge_pump_2/in3 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 35.68658f
C614 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C615 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C616 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C617 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C618 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C619 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C620 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C621 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C622 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C623 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C624 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C625 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C626 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C627 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C628 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C629 CP2_5_stage_0/charge_pump_0/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.390842f
C630 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C631 CP2_5_stage_0/charge_pump_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 84.016754f
C632 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C633 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C634 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C635 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C636 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C637 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C638 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C639 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C640 CP2_5_stage_0/charge_pump_0/g1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.668617f
C641 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.79532f
C642 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C643 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C644 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C645 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C646 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C647 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C648 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.234749f
C649 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C650 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C651 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C652 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C653 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C654 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C655 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C656 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C657 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C658 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C659 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C660 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C661 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C662 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C663 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C664 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/out1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.075895f
C665 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C666 CP2_5_stage_1/charge_pump_reverse_1/clock_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 90.940094f
C667 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C668 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C669 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C670 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C671 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C672 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C673 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C674 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C675 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C676 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C677 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C678 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C679 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C680 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C681 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C682 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C683 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C684 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C685 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C686 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C687 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C688 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C689 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C690 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/out2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.860609f
C691 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C692 CP2_5_stage_1/charge_pump_reverse_1/clock_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 84.53275f
C693 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C694 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C695 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C696 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C697 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C698 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C699 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C700 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C701 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.425359f
C702 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.79532f
C703 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C704 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C705 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C706 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C707 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C708 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C709 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.234749f
C710 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C711 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C712 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C713 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C714 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C715 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C716 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C717 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C718 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C719 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C720 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C721 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C722 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C723 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C724 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C725 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/out1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.076454f
C726 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C727 CP2_5_stage_1/charge_pump_reverse_0/clock_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 90.94089f
C728 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C729 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C730 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C731 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C732 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C733 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C734 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C735 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C736 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C737 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C738 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C739 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C740 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C741 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C742 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C743 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C744 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C745 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C746 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C747 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C748 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C749 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C750 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C751 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/out2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.861251f
C752 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C753 CP2_5_stage_1/charge_pump_reverse_0/clock_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 84.53365f
C754 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C755 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C756 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C757 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C758 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C759 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C760 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C761 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C762 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.425359f
C763 CP2_5_stage_1/buffer_digital_6/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 10.263865f
C764 CP2_5_stage_1/buffer_digital_2/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.585812f
C765 CP2_5_stage_1/charge_pump_2/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.96237f
C766 CP2_5_stage_1/charge_pump_2/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C767 CP2_5_stage_1/charge_pump_2/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C768 CP2_5_stage_1/charge_pump_2/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C769 CP2_5_stage_1/charge_pump_2/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C770 CP2_5_stage_1/charge_pump_2/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C771 CP2_5_stage_1/buffer_digital_7/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 17.893332f
C772 CP2_5_stage_1/charge_pump_2/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C773 CP2_5_stage_1/charge_pump_2/g2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.43748f
C774 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C775 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C776 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C777 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C778 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C779 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C780 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C781 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C782 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C783 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C784 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C785 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C786 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C787 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C788 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C789 CP2_5_stage_1/charge_pump_2/in1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 49.778893f
C790 CP2_5_stage_1/charge_pump_2/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.031953f
C791 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C792 CP2_5_stage_1/charge_pump_2/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 82.29622f
C793 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C794 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C795 CP2_5_stage_1/charge_pump_2/in8 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 57.29606f
C796 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C797 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C798 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C799 CP2_5_stage_1/charge_pump_2/in7 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 50.83537f
C800 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C801 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C802 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C803 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C804 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C805 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C806 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C807 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C808 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C809 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C810 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C811 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C812 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C813 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C814 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C815 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C816 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C817 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C818 CP2_5_stage_1/charge_pump_2/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.390842f
C819 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C820 CP2_5_stage_1/charge_pump_2/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 83.97966f
C821 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C822 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C823 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C824 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C825 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C826 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C827 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C828 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C829 CP2_5_stage_1/charge_pump_2/g1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.634558f
C830 CP2_5_stage_1/buffer_digital_1/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.342446f
C831 CP2_5_stage_1/charge_pump_1/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.96237f
C832 CP2_5_stage_1/charge_pump_1/out CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 3.305988f
C833 CP2_5_stage_1/charge_pump_1/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C834 CP2_5_stage_1/charge_pump_1/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C835 CP2_5_stage_1/charge_pump_1/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C836 CP2_5_stage_1/charge_pump_1/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C837 CP2_5_stage_1/charge_pump_1/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C838 CP2_5_stage_1/buffer_digital_4/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.588428f
C839 CP2_5_stage_1/charge_pump_1/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C840 CP2_5_stage_1/charge_pump_1/g2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.43748f
C841 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C842 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C843 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C844 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C845 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C846 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C847 CP2_5_stage_1/charge_pump_2/in4 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 32.558914f
C848 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C849 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C850 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C851 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C852 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C853 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C854 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C855 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C856 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C857 CP2_5_stage_1/charge_pump_1/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.031953f
C858 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C859 CP2_5_stage_1/charge_pump_1/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 82.29622f
C860 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C861 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C862 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C863 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C864 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C865 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C866 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C867 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C868 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C869 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C870 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C871 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C872 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C873 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C874 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C875 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C876 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C877 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C878 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C879 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C880 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C881 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C882 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C883 CP2_5_stage_1/charge_pump_1/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.390842f
C884 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C885 CP2_5_stage_1/charge_pump_1/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 83.97966f
C886 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C887 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C888 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C889 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C890 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C891 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C892 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C893 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C894 CP2_5_stage_1/charge_pump_1/g1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.634558f
C895 CP2_5_stage_1/charge_pump_0/vin CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 3.426366f
C896 CP2_5_stage_1/charge_pump_0/vs CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 18.96202f
C897 CP2_5_stage_1/charge_pump_0/clock_0/a_2432_n962# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 8.68424f **FLOATING
C898 CP2_5_stage_1/charge_pump_0/clock_0/a_2020_n482# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.56615f **FLOATING
C899 CP2_5_stage_1/charge_pump_0/clock_0/a_344_102# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.809951f
C900 CP2_5_stage_1/charge_pump_0/clock_0/a_2402_572# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.172722f
C901 CP2_5_stage_1/charge_pump_0/clock_0/a_344_n986# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.381627f
C902 CP2_5_stage_1/buffer_digital_0/i CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 0.107092p
C903 CP2_5_stage_1/charge_pump_0/clock_0/a_3246_118# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.834443f
C904 CP2_5_stage_1/charge_pump_0/g2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.43748f
C905 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C906 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C907 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C908 CP2_5_stage_1/charge_pump_2/in5 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 33.069042f
C909 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C910 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C911 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C912 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C913 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C914 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C915 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C916 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C917 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C918 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C919 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C920 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C921 CP2_5_stage_1/charge_pump_0/input1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 15.031953f
C922 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C923 CP2_5_stage_1/charge_pump_0/clk CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 82.25907f
C924 CP1_5_stage_0/charge_pump1_2/vdd CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 6.971405p
C925 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C926 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C927 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C928 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C929 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C930 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C931 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C932 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C933 CP2_5_stage_1/charge_pump_2/in6 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 44.152824f
C934 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C935 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C936 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C937 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C938 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C939 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C940 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C941 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C942 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C943 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C944 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C945 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C946 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C947 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C948 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C949 CP2_5_stage_1/charge_pump_0/input2 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 14.390842f
C950 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C951 CP2_5_stage_1/charge_pump_0/clkb CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 83.97966f
C952 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C953 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C954 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C955 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C956 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C957 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.337696f
C958 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 9.978376f
C959 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.581652f
C960 CP2_5_stage_1/charge_pump_0/g1 CP2_5_stage_0/charge_pump_2/nmos_diode2_0/VSUBS 2.634558f
.ends

