magic
tech sky130A
magscale 1 2
timestamp 1699221170
<< metal1 >>
rect 104638 28312 105070 28318
rect 104638 28248 104680 28312
rect 105054 28248 105070 28312
rect 104638 28246 104774 28248
rect 104922 28246 105070 28248
rect 104638 28234 105070 28246
rect 104744 28232 104950 28234
rect -3758 26622 -3492 26666
rect -3780 26540 -3492 26622
rect -3780 25918 -3708 26540
rect -3538 25918 -3492 26540
rect -3780 25872 -3492 25918
rect -3780 -18670 -3604 25872
rect -3790 -18790 -3604 -18670
rect -3790 -19380 -3768 -18790
rect -3636 -19380 -3604 -18790
rect -3790 -19452 -3604 -19380
rect -3780 -50248 -3604 -19452
rect -3454 24396 -3244 24525
rect -3454 23774 -3432 24396
rect -3262 23774 -3244 24396
rect -3454 -16812 -3244 23774
rect -3454 -17402 -3428 -16812
rect -3296 -17402 -3244 -16812
rect -3454 -48132 -3244 -17402
rect -2934 22322 -2682 22414
rect -2934 21700 -2884 22322
rect -2714 21700 -2682 22322
rect -2934 -14686 -2682 21700
rect -2934 -15276 -2894 -14686
rect -2762 -15276 -2682 -14686
rect -2934 -46138 -2682 -15276
rect -2454 20256 -2202 20340
rect -2454 19634 -2410 20256
rect -2240 19634 -2202 20256
rect -2454 -12634 -2202 19634
rect -2454 -13224 -2396 -12634
rect -2264 -13224 -2202 -12634
rect -2454 -44068 -2202 -13224
rect -1942 18154 -1690 18260
rect -1942 17532 -1914 18154
rect -1744 17532 -1690 18154
rect -1942 -10482 -1690 17532
rect -1942 -11066 -1936 -10482
rect -1762 -10694 -1690 -10482
rect -1504 16102 -1252 16128
rect -1504 15480 -1458 16102
rect -1288 15480 -1252 16102
rect -1504 -8532 -1252 15480
rect -1066 13920 -800 14038
rect -1066 13298 -1026 13920
rect -856 13298 -800 13920
rect -1066 13244 -800 13298
rect -1052 -6306 -800 13244
rect -440 11850 -188 11862
rect -460 11782 -124 11850
rect -460 11160 -350 11782
rect -180 11160 -124 11782
rect -460 11082 -124 11160
rect -1066 -6406 -800 -6306
rect -1066 -6990 -1016 -6406
rect -842 -6520 -800 -6406
rect -440 -4428 -188 11082
rect 94628 -348 95574 -338
rect 94626 -374 95574 -348
rect 94626 -486 94694 -374
rect 95496 -486 95574 -374
rect 94626 -528 95574 -486
rect 24666 -2758 24986 -2712
rect 24666 -2934 24702 -2758
rect 24928 -2934 24986 -2758
rect 26684 -2787 26696 -2651
rect 47710 -2658 48120 -2651
rect 47710 -2734 48286 -2658
rect 47710 -2787 48124 -2734
rect 24666 -2952 24986 -2934
rect -440 -5034 -382 -4428
rect -262 -5034 -188 -4428
rect -842 -6990 -778 -6520
rect -1066 -7100 -778 -6990
rect -1504 -9116 -1462 -8532
rect -1288 -9116 -1252 -8532
rect -1762 -11066 -1684 -10694
rect -1942 -41992 -1684 -11066
rect -1504 -39904 -1252 -9116
rect -1052 -37712 -778 -7100
rect -440 -35698 -188 -5034
rect 22331 -21160 24560 -21030
rect 24750 -21656 24886 -2952
rect 48084 -3376 48124 -2787
rect 48242 -3376 48286 -2734
rect 94626 -2753 94762 -528
rect 48084 -3426 48286 -3376
rect 104762 -3469 104920 28232
rect 71703 -20442 71833 -20435
rect 71606 -20532 71932 -20442
rect 71606 -21006 71690 -20532
rect 70369 -21086 71690 -21006
rect 71866 -21086 71932 -20532
rect 70369 -21136 71932 -21086
rect 71606 -21138 71932 -21136
rect 24706 -21732 24890 -21656
rect 24706 -22182 24734 -21732
rect 24838 -22182 24890 -21732
rect 24706 -22228 24890 -22182
rect 24750 -22232 24886 -22228
rect 24340 -31862 24810 -31782
rect 24340 -32064 24390 -31862
rect 24754 -31956 24810 -31862
rect 24754 -32064 24830 -31956
rect 24340 -32084 24830 -32064
rect 24340 -32114 24810 -32084
rect 24350 -35203 24478 -32114
rect 72400 -34373 72784 -34372
rect 72400 -34450 73316 -34373
rect 72400 -35080 72502 -34450
rect 72720 -34509 73316 -34450
rect 72720 -35080 72784 -34509
rect 72400 -35162 72784 -35080
rect -440 -36180 -382 -35698
rect -240 -36180 -188 -35698
rect -440 -36262 -188 -36180
rect -250 -36315 -196 -36262
rect -1058 -37778 -778 -37712
rect -1058 -38260 -998 -37778
rect -856 -38260 -778 -37778
rect -1058 -38366 -778 -38260
rect -850 -38368 -778 -38366
rect -1504 -40386 -1436 -39904
rect -1294 -40386 -1252 -39904
rect -1504 -40440 -1252 -40386
rect -1332 -40462 -1268 -40440
rect -1942 -42474 -1854 -41992
rect -1712 -42474 -1684 -41992
rect -1942 -42549 -1684 -42474
rect -1942 -42552 -1690 -42549
rect -2454 -44550 -2388 -44068
rect -2246 -44550 -2202 -44068
rect -2454 -44624 -2202 -44550
rect -2270 -44639 -2224 -44624
rect -2934 -46620 -2894 -46138
rect -2752 -46620 -2682 -46138
rect -2934 -46718 -2682 -46620
rect -3454 -48230 -3196 -48132
rect -3454 -48712 -3394 -48230
rect -3252 -48712 -3196 -48230
rect -3454 -48786 -3196 -48712
rect -3454 -48790 -3244 -48786
rect -3306 -48899 -3244 -48790
rect -3796 -50356 -3538 -50248
rect -3796 -50838 -3744 -50356
rect -3602 -50838 -3538 -50356
rect -3796 -50902 -3538 -50838
rect -3780 -50918 -3604 -50902
rect 48961 -52224 49242 -52162
rect 48961 -52818 49002 -52224
rect 49184 -52728 49242 -52224
rect 95919 -52276 96160 -52178
rect 49184 -52818 51491 -52728
rect 48961 -52858 51491 -52818
rect 95919 -52828 95992 -52276
rect 96120 -52752 96160 -52276
rect 96120 -52828 98511 -52752
rect 95919 -52882 98511 -52828
<< via1 >>
rect 104680 28248 105054 28312
rect 104774 28246 104922 28248
rect -3708 25918 -3538 26540
rect -3768 -19380 -3636 -18790
rect -3432 23774 -3262 24396
rect -3428 -17402 -3296 -16812
rect -2884 21700 -2714 22322
rect -2894 -15276 -2762 -14686
rect -2410 19634 -2240 20256
rect -2396 -13224 -2264 -12634
rect -1914 17532 -1744 18154
rect -1936 -11066 -1762 -10482
rect -1458 15480 -1288 16102
rect -1026 13298 -856 13920
rect -350 11160 -180 11782
rect -1016 -6990 -842 -6406
rect 94694 -486 95496 -374
rect 24702 -2934 24928 -2758
rect -382 -5034 -262 -4428
rect -1462 -9116 -1288 -8532
rect 48124 -3376 48242 -2734
rect 71690 -21086 71866 -20532
rect 24734 -22182 24838 -21732
rect 24390 -32064 24754 -31862
rect 72502 -35080 72720 -34450
rect -382 -36180 -240 -35698
rect -998 -38260 -856 -37778
rect -1436 -40386 -1294 -39904
rect -1854 -42474 -1712 -41992
rect -2388 -44550 -2246 -44068
rect -2894 -46620 -2752 -46138
rect -3394 -48712 -3252 -48230
rect -3744 -50838 -3602 -50356
rect 49002 -52818 49184 -52224
rect 95992 -52828 96120 -52276
<< metal2 >>
rect -3758 26628 -3492 26666
rect -3767 26582 2969 26628
rect -3758 26540 -3492 26582
rect -3758 25918 -3708 26540
rect -3538 25918 -3492 26540
rect -3758 25872 -3492 25918
rect -3459 24500 2939 24522
rect -3482 24476 2939 24500
rect -3482 24396 -3216 24476
rect -3482 23774 -3432 24396
rect -3262 23774 -3216 24396
rect -3482 23706 -3216 23774
rect -2926 22428 -2660 22430
rect -2931 22382 2939 22428
rect -2926 22322 -2660 22382
rect -2926 21700 -2884 22322
rect -2714 21700 -2660 22322
rect -2926 21636 -2660 21700
rect -2456 20334 -2190 20346
rect -2456 20288 2937 20334
rect -2456 20256 -2190 20288
rect -2456 19634 -2410 20256
rect -2240 19634 -2190 20256
rect -2456 19552 -2190 19634
rect -1941 18238 2919 18240
rect -1954 18194 2919 18238
rect -1954 18154 -1688 18194
rect -1954 17532 -1914 18154
rect -1744 17532 -1688 18154
rect -1954 17444 -1688 17532
rect -1494 16146 -1228 16178
rect -1537 16102 2929 16146
rect -1537 16100 -1458 16102
rect -1494 15480 -1458 16100
rect -1288 16100 2929 16102
rect -1288 15480 -1228 16100
rect -1494 15384 -1228 15480
rect -1067 14006 2931 14052
rect -1066 13920 -800 14006
rect -1066 13298 -1026 13920
rect -856 13298 -800 13920
rect -1066 13244 -800 13298
rect -414 11864 -148 11876
rect -463 11810 3028 11864
rect -414 11782 -148 11810
rect -414 11160 -350 11782
rect -180 11160 -148 11782
rect -414 11082 -148 11160
rect 127438 10042 132222 10126
rect 94628 -374 123398 -338
rect 94628 -486 94694 -374
rect 95496 -402 123398 -374
rect 95496 -486 95574 -402
rect 94628 -528 95574 -486
rect 48084 -2734 48286 -2658
rect 48084 -3367 48124 -2734
rect 48082 -3376 48124 -3367
rect 48242 -3367 48286 -2734
rect 123334 -3341 123398 -402
rect 132138 -3341 132222 10042
rect 48242 -3376 50406 -3367
rect 48082 -3431 50406 -3376
rect 114708 -3405 132254 -3341
rect 132138 -3416 132222 -3405
rect -450 -4428 -184 -4318
rect -450 -5034 -382 -4428
rect -262 -4554 -184 -4428
rect -262 -4602 2955 -4554
rect -262 -4609 681 -4602
rect -262 -5034 -184 -4609
rect -450 -5112 -184 -5034
rect -1066 -6406 -800 -6306
rect -1066 -6990 -1016 -6406
rect -842 -6633 -800 -6406
rect -842 -6681 2976 -6633
rect -842 -6990 -800 -6681
rect -1066 -7100 -800 -6990
rect -1500 -8532 -1234 -8394
rect -1500 -8727 -1462 -8532
rect -1518 -8775 -1462 -8727
rect -1500 -9116 -1462 -8775
rect -1288 -8727 -1234 -8532
rect -1288 -8775 2974 -8727
rect -1288 -9116 -1234 -8775
rect -1500 -9188 -1234 -9116
rect -1968 -10482 -1702 -10386
rect -1968 -10817 -1936 -10482
rect -2434 -10865 -1936 -10817
rect -1968 -11066 -1936 -10865
rect -1762 -10817 -1702 -10482
rect -1762 -10865 3064 -10817
rect -1762 -11066 -1702 -10865
rect -1968 -11180 -1702 -11066
rect -2460 -12634 -2226 -12516
rect -2460 -12918 -2396 -12634
rect -2472 -12966 -2396 -12918
rect -2460 -13224 -2396 -12966
rect -2264 -12918 -2226 -12634
rect -2264 -12966 3043 -12918
rect -2264 -13224 -2226 -12966
rect -2460 -13298 -2226 -13224
rect -2944 -14686 -2710 -14554
rect -2944 -15276 -2894 -14686
rect -2762 -14997 -2710 -14686
rect -2762 -15045 3058 -14997
rect -2762 -15276 -2710 -15045
rect -2944 -15336 -2710 -15276
rect -3446 -16812 -3266 -16692
rect -3446 -17402 -3428 -16812
rect -3296 -17091 -3266 -16812
rect -3296 -17139 3062 -17091
rect -3296 -17402 -3266 -17139
rect -3446 -17474 -3266 -17402
rect -3790 -18790 -3616 -18670
rect -3790 -19380 -3768 -18790
rect -3636 -19177 -3616 -18790
rect -3636 -19225 3056 -19177
rect -3636 -19380 -3616 -19225
rect -3790 -19452 -3616 -19380
rect 71685 -20442 73831 -20435
rect 71606 -20532 73831 -20442
rect 9894 -35210 10134 -21017
rect 71606 -21086 71690 -20532
rect 71866 -20549 73831 -20532
rect 71866 -21086 71932 -20549
rect 71606 -21138 71932 -21086
rect 24706 -21732 24890 -21656
rect 24706 -22182 24734 -21732
rect 24838 -22182 24890 -21732
rect 24706 -22228 24890 -22182
rect 24709 -31782 24823 -22228
rect 24340 -31862 24823 -31782
rect 24340 -32064 24390 -31862
rect 24754 -32064 24823 -31862
rect 24340 -32083 24823 -32064
rect 24340 -32114 24810 -32083
rect 72342 -34450 72810 -34378
rect 72342 -35080 72502 -34450
rect 72720 -35080 72810 -34450
rect 72342 -35089 72810 -35080
rect 71268 -35153 72810 -35089
rect -442 -35698 -184 -35606
rect -442 -36180 -382 -35698
rect -240 -36180 -184 -35698
rect -442 -36225 -184 -36180
rect -442 -36260 3662 -36225
rect -254 -36273 3662 -36260
rect -1058 -37778 -800 -37712
rect -1058 -38260 -998 -37778
rect -856 -38260 -800 -37778
rect -1058 -38311 -800 -38260
rect -1058 -38359 3674 -38311
rect -1058 -38366 -800 -38359
rect -1514 -39904 -1256 -39810
rect -1514 -40386 -1436 -39904
rect -1294 -40386 -1256 -39904
rect -1514 -40405 -1256 -40386
rect -1514 -40453 3654 -40405
rect -1514 -40464 -1256 -40453
rect -1918 -41992 -1660 -41884
rect -1918 -42474 -1854 -41992
rect -1712 -42474 -1660 -41992
rect -1918 -42495 -1660 -42474
rect -1918 -42538 3738 -42495
rect -1784 -42543 3738 -42538
rect -2452 -44068 -2194 -43978
rect -2452 -44550 -2388 -44068
rect -2246 -44550 -2194 -44068
rect -2452 -44593 -2194 -44550
rect -2452 -44632 3730 -44593
rect -2260 -44641 3730 -44632
rect -2958 -46138 -2700 -46076
rect -2958 -46620 -2894 -46138
rect -2752 -46620 -2700 -46138
rect -2958 -46675 -2700 -46620
rect -2958 -46723 3718 -46675
rect -2958 -46730 -2700 -46723
rect -3454 -48230 -3196 -48132
rect -3454 -48712 -3394 -48230
rect -3252 -48712 -3196 -48230
rect -3454 -48769 -3196 -48712
rect -3454 -48786 3720 -48769
rect -3302 -48817 3720 -48786
rect -3796 -50356 -3538 -50248
rect -3796 -50838 -3744 -50356
rect -3602 -50838 -3538 -50356
rect -3796 -50855 -3538 -50838
rect -3796 -50902 3728 -50855
rect -3774 -50903 3728 -50902
rect 46993 -52162 49109 -52157
rect 46993 -52224 49242 -52162
rect 95919 -52191 96160 -52178
rect 46993 -52271 49002 -52224
rect 48961 -52818 49002 -52271
rect 49184 -52818 49242 -52224
rect 93843 -52276 96160 -52191
rect 93843 -52305 95992 -52276
rect 48961 -52858 49242 -52818
rect 95919 -52828 95992 -52305
rect 96120 -52828 96160 -52276
rect 95919 -52882 96160 -52828
<< metal3 >>
rect 412 1112 804 1262
rect 379 734 7415 1112
rect 412 -32254 804 734
rect 118478 -30419 118870 -30354
rect 113438 -30811 119110 -30419
rect 118478 -31476 118870 -30811
rect 29784 -31568 60480 -31476
rect 61948 -31538 107514 -31476
rect 108948 -31538 118870 -31476
rect 61948 -31568 118870 -31538
rect 29784 -31868 118870 -31568
rect 29784 -32254 30176 -31868
rect 412 -32646 30176 -32254
rect 412 -62141 804 -32646
rect 412 -62533 5806 -62141
rect 117768 -62601 119110 -62209
<< metal4 >>
rect 118772 -4699 119470 1755
rect 118772 -35777 119470 -29431
<< metal5 >>
rect 117867 -2420 118525 703
rect 119748 -37415 120466 -29963
use cp1_buffer_5stage  cp1_buffer_5stage_0
timestamp 1699130246
transform 1 0 1331 0 1 130
box -1331 -130 130524 30508
use cp2_buffer_5stage  cp2_buffer_5stage_0
timestamp 1699177610
transform -1 0 95205 0 1 -31824
box -25261 108 95113 31581
use cp2_buffer_5stage  cp2_buffer_5stage_1
timestamp 1699177610
transform 1 0 25637 0 1 -63546
box -25261 108 95113 31581
<< end >>
