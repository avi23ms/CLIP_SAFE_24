magic
tech sky130A
magscale 1 2
timestamp 1699177610
<< dnwell >>
rect 12148 -412 12324 -348
<< nwell >>
rect 22756 16112 23104 16396
rect 1550 8230 1848 8398
<< psubdiff >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
<< nsubdiff >>
rect 12178 17270 12374 17296
rect 12178 17166 12210 17270
rect 12338 17166 12374 17270
rect 12178 17134 12374 17166
rect 22804 16354 22876 16356
rect 22794 16330 22878 16354
rect 22794 16190 22818 16330
rect 22854 16192 22878 16330
rect 22852 16190 22878 16192
rect 22794 16164 22878 16190
rect 1662 8334 1794 8360
rect 1662 8294 1692 8334
rect 1758 8294 1794 8334
rect 1662 8270 1794 8294
rect 12180 684 12366 716
rect 12180 578 12216 684
rect 12334 578 12366 684
rect 12180 554 12366 578
<< psubdiffcont >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
<< nsubdiffcont >>
rect 12210 17166 12338 17270
rect 22818 16192 22854 16330
rect 22818 16190 22852 16192
rect 1692 8294 1758 8334
rect 12216 578 12334 684
<< poly >>
rect 1442 16632 1516 16694
rect 1424 16602 1516 16632
rect 1442 16440 1516 16602
rect 1422 16410 1516 16440
rect 1442 16248 1516 16410
rect 1422 16218 1516 16248
rect 1442 16056 1516 16218
rect 23136 16296 23224 16652
rect 23106 16266 23224 16296
rect 23136 16104 23224 16266
rect 23106 16074 23224 16104
rect 1418 16026 1516 16056
rect 1442 15864 1516 16026
rect 23136 15912 23224 16074
rect 23106 15882 23224 15912
rect 1422 15834 1516 15864
rect 1442 15672 1516 15834
rect 23136 15720 23224 15882
rect 23104 15690 23224 15720
rect 1420 15642 1516 15672
rect 1442 15480 1516 15642
rect 23136 15528 23224 15690
rect 23104 15498 23224 15528
rect 1418 15450 1516 15480
rect 1442 15288 1516 15450
rect 23136 15336 23224 15498
rect 23104 15306 23224 15336
rect 1422 15258 1516 15288
rect 1442 15096 1516 15258
rect 23136 15144 23224 15306
rect 23106 15114 23224 15144
rect 1422 15066 1516 15096
rect 1442 14904 1516 15066
rect 23136 14952 23224 15114
rect 23106 14922 23224 14952
rect 1422 14874 1516 14904
rect 1442 14712 1516 14874
rect 23136 14760 23224 14922
rect 23104 14730 23224 14760
rect 1422 14682 1516 14712
rect 1442 14520 1516 14682
rect 23136 14568 23224 14730
rect 23106 14538 23224 14568
rect 1420 14490 1516 14520
rect 1442 14328 1516 14490
rect 23136 14376 23224 14538
rect 23106 14346 23224 14376
rect 1424 14298 1516 14328
rect 1442 14136 1516 14298
rect 23136 14184 23224 14346
rect 23102 14154 23224 14184
rect 1420 14106 1516 14136
rect 1442 13944 1516 14106
rect 23136 13992 23224 14154
rect 23102 13962 23224 13992
rect 1422 13914 1516 13944
rect 1442 13752 1516 13914
rect 23136 13800 23224 13962
rect 23104 13770 23224 13800
rect 1420 13722 1516 13752
rect 1442 13560 1516 13722
rect 23136 13608 23224 13770
rect 23108 13578 23224 13608
rect 1422 13530 1516 13560
rect 1442 13368 1516 13530
rect 23136 13416 23224 13578
rect 23100 13386 23224 13416
rect 1422 13338 1516 13368
rect 1442 13176 1516 13338
rect 23136 13224 23224 13386
rect 23104 13194 23224 13224
rect 1418 13146 1516 13176
rect 1442 12984 1516 13146
rect 23136 13032 23224 13194
rect 23102 13002 23224 13032
rect 1416 12954 1516 12984
rect 1442 12792 1516 12954
rect 23136 12840 23224 13002
rect 23104 12810 23224 12840
rect 1422 12762 1516 12792
rect 1442 12600 1516 12762
rect 23136 12648 23224 12810
rect 23104 12618 23224 12648
rect 1422 12570 1516 12600
rect 1442 12408 1516 12570
rect 23136 12456 23224 12618
rect 23104 12426 23224 12456
rect 1418 12378 1516 12408
rect 1442 12216 1516 12378
rect 23136 12264 23224 12426
rect 23100 12234 23224 12264
rect 1420 12186 1516 12216
rect 1442 12024 1516 12186
rect 23136 12072 23224 12234
rect 23100 12042 23224 12072
rect 1418 11994 1516 12024
rect 1442 11832 1516 11994
rect 23136 11880 23224 12042
rect 23106 11850 23224 11880
rect 1420 11802 1516 11832
rect 1442 11640 1516 11802
rect 23136 11688 23224 11850
rect 23104 11658 23224 11688
rect 1418 11610 1516 11640
rect 1442 11448 1516 11610
rect 23136 11496 23224 11658
rect 23104 11466 23224 11496
rect 1420 11418 1516 11448
rect 1442 11256 1516 11418
rect 23136 11304 23224 11466
rect 23104 11274 23224 11304
rect 1418 11226 1516 11256
rect 1442 11064 1516 11226
rect 23136 11112 23224 11274
rect 23098 11082 23224 11112
rect 1420 11034 1516 11064
rect 1442 10872 1516 11034
rect 23136 10920 23224 11082
rect 23100 10890 23224 10920
rect 1420 10842 1516 10872
rect 1442 10680 1516 10842
rect 23136 10728 23224 10890
rect 23100 10698 23224 10728
rect 1424 10650 1516 10680
rect 1442 10488 1516 10650
rect 23136 10536 23224 10698
rect 23102 10506 23224 10536
rect 1424 10458 1516 10488
rect 1442 10296 1516 10458
rect 23136 10344 23224 10506
rect 23098 10314 23224 10344
rect 1422 10266 1516 10296
rect 1442 10104 1516 10266
rect 23136 10152 23224 10314
rect 23102 10122 23224 10152
rect 1424 10074 1516 10104
rect 1442 9912 1516 10074
rect 23136 9960 23224 10122
rect 23102 9930 23224 9960
rect 1424 9882 1516 9912
rect 1442 9720 1516 9882
rect 23136 9768 23224 9930
rect 23104 9738 23224 9768
rect 1424 9690 1516 9720
rect 1442 9528 1516 9690
rect 23136 9576 23224 9738
rect 23102 9546 23224 9576
rect 1424 9498 1516 9528
rect 1442 9336 1516 9498
rect 23136 9384 23224 9546
rect 23098 9354 23224 9384
rect 1422 9306 1516 9336
rect 1442 9144 1516 9306
rect 23136 9192 23224 9354
rect 23102 9162 23224 9192
rect 1416 9114 1516 9144
rect 1442 8912 1516 9114
rect 23136 9000 23224 9162
rect 23096 8970 23224 9000
rect 23136 8808 23224 8970
rect 23092 8778 23224 8808
rect 23136 8554 23224 8778
rect 1262 8196 1384 8416
rect 1262 8166 1428 8196
rect 1262 8004 1384 8166
rect 1262 7974 1438 8004
rect 1262 7812 1384 7974
rect 1262 7782 1428 7812
rect 1262 7620 1384 7782
rect 23000 7758 23152 7934
rect 23000 7728 23194 7758
rect 1262 7590 1436 7620
rect 1262 7428 1384 7590
rect 23000 7566 23152 7728
rect 23000 7536 23196 7566
rect 1262 7398 1436 7428
rect 1262 7236 1384 7398
rect 23000 7374 23152 7536
rect 23000 7344 23194 7374
rect 1262 7206 1432 7236
rect 1262 7044 1384 7206
rect 23000 7182 23152 7344
rect 23000 7152 23192 7182
rect 1262 7014 1432 7044
rect 1262 6852 1384 7014
rect 23000 6990 23152 7152
rect 23000 6960 23198 6990
rect 1262 6822 1440 6852
rect 1262 6660 1384 6822
rect 23000 6798 23152 6960
rect 23000 6768 23204 6798
rect 1262 6630 1430 6660
rect 1262 6468 1384 6630
rect 23000 6606 23152 6768
rect 23000 6576 23198 6606
rect 1262 6438 1438 6468
rect 1262 6276 1384 6438
rect 23000 6414 23152 6576
rect 23000 6384 23200 6414
rect 1262 6246 1432 6276
rect 1262 6084 1384 6246
rect 23000 6222 23152 6384
rect 23000 6192 23206 6222
rect 1262 6054 1440 6084
rect 1262 5892 1384 6054
rect 23000 6030 23152 6192
rect 23000 6000 23196 6030
rect 1262 5862 1440 5892
rect 1262 5700 1384 5862
rect 23000 5838 23152 6000
rect 23000 5808 23200 5838
rect 1262 5670 1436 5700
rect 1262 5508 1384 5670
rect 23000 5646 23152 5808
rect 23000 5616 23198 5646
rect 1262 5478 1440 5508
rect 1262 5316 1384 5478
rect 23000 5454 23152 5616
rect 23000 5424 23200 5454
rect 1262 5286 1434 5316
rect 1262 5124 1384 5286
rect 23000 5262 23152 5424
rect 23000 5232 23204 5262
rect 1262 5094 1440 5124
rect 1262 4932 1384 5094
rect 23000 5070 23152 5232
rect 23000 5040 23200 5070
rect 1262 4902 1440 4932
rect 1262 4740 1384 4902
rect 23000 4878 23152 5040
rect 23000 4848 23208 4878
rect 1262 4710 1430 4740
rect 1262 4548 1384 4710
rect 23000 4686 23152 4848
rect 23000 4656 23198 4686
rect 1262 4518 1426 4548
rect 1262 4356 1384 4518
rect 23000 4494 23152 4656
rect 23000 4464 23194 4494
rect 1262 4326 1436 4356
rect 1262 4164 1384 4326
rect 23000 4302 23152 4464
rect 23000 4272 23198 4302
rect 1262 4134 1442 4164
rect 1262 3972 1384 4134
rect 23000 4110 23152 4272
rect 23000 4080 23198 4110
rect 1262 3942 1444 3972
rect 1262 3780 1384 3942
rect 23000 3918 23152 4080
rect 23000 3888 23196 3918
rect 1262 3750 1440 3780
rect 1262 3588 1384 3750
rect 23000 3726 23152 3888
rect 23000 3696 23194 3726
rect 1262 3558 1440 3588
rect 1262 3396 1384 3558
rect 23000 3534 23152 3696
rect 23000 3504 23200 3534
rect 1262 3366 1438 3396
rect 1262 3204 1384 3366
rect 23000 3342 23152 3504
rect 23000 3312 23196 3342
rect 1262 3174 1430 3204
rect 1262 3012 1384 3174
rect 23000 3150 23152 3312
rect 23000 3120 23198 3150
rect 1262 2982 1438 3012
rect 1262 2820 1384 2982
rect 23000 2958 23152 3120
rect 23000 2928 23204 2958
rect 1262 2790 1440 2820
rect 1262 2628 1384 2790
rect 23000 2766 23152 2928
rect 23000 2736 23196 2766
rect 1262 2598 1434 2628
rect 1262 2436 1384 2598
rect 23000 2574 23152 2736
rect 23000 2544 23198 2574
rect 1262 2406 1434 2436
rect 1262 2244 1384 2406
rect 23000 2382 23152 2544
rect 23000 2352 23196 2382
rect 1262 2214 1440 2244
rect 1262 2052 1384 2214
rect 23000 2190 23152 2352
rect 23000 2160 23194 2190
rect 1262 2022 1442 2052
rect 1262 1860 1384 2022
rect 23000 1998 23152 2160
rect 23000 1968 23192 1998
rect 1262 1830 1440 1860
rect 1262 1668 1384 1830
rect 23000 1806 23152 1968
rect 23000 1776 23194 1806
rect 1262 1638 1438 1668
rect 1262 1476 1384 1638
rect 23000 1614 23152 1776
rect 23000 1584 23198 1614
rect 1262 1446 1440 1476
rect 1262 1284 1384 1446
rect 23000 1422 23152 1584
rect 23000 1392 23198 1422
rect 1262 1254 1438 1284
rect 1262 1092 1384 1254
rect 23000 1230 23152 1392
rect 23000 1200 23206 1230
rect 1262 1062 1432 1092
rect 1262 900 1384 1062
rect 23000 1038 23152 1200
rect 23000 1008 23196 1038
rect 1262 870 1442 900
rect 1262 708 1384 870
rect 23000 846 23152 1008
rect 23000 816 23200 846
rect 1262 678 1444 708
rect 1262 558 1384 678
rect 23000 654 23152 816
rect 23000 624 23196 654
rect 23000 462 23152 624
rect 23000 432 23202 462
rect 23000 270 23152 432
rect 23000 240 23198 270
rect 23000 208 23152 240
<< locali >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
rect 12178 17270 12374 17296
rect 12178 17166 12210 17270
rect 12338 17166 12374 17270
rect 12178 17134 12374 17166
rect 1494 16694 1932 16696
rect 1442 16576 1932 16694
rect 1442 8950 1692 16576
rect 1838 8950 1932 16576
rect 23136 16412 23714 16674
rect 22804 16354 22876 16356
rect 22794 16330 22878 16354
rect 22794 16190 22818 16330
rect 22854 16192 22878 16330
rect 22852 16190 22878 16192
rect 22794 16164 22878 16190
rect 1442 8912 1932 8950
rect 1494 8908 1932 8912
rect 894 8416 1314 8806
rect 23136 8756 23332 16412
rect 23638 8756 23714 16412
rect 23136 8554 23714 8756
rect 894 8338 1388 8416
rect 894 696 1006 8338
rect 1214 696 1388 8338
rect 1662 8334 1794 8360
rect 1662 8294 1692 8334
rect 1758 8294 1794 8334
rect 1662 8270 1794 8294
rect 22746 7934 23096 7936
rect 22614 7930 23096 7934
rect 22614 7792 23152 7930
rect 894 584 1388 696
rect 1096 552 1388 584
rect 12182 684 12368 714
rect 12182 578 12216 684
rect 12334 578 12368 684
rect 12182 552 12368 578
rect 22614 278 22698 7792
rect 22980 278 23152 7792
rect 22614 114 23152 278
rect 22614 110 23004 114
rect 13076 48 13132 52
rect 13076 -216 13132 -214
<< viali >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 12210 17166 12338 17270
rect 1692 8950 1838 16576
rect 22818 16190 22852 16330
rect 23332 8756 23638 16412
rect 1006 696 1214 8338
rect 1692 8294 1758 8334
rect 12216 578 12334 684
rect 22698 278 22980 7792
rect 13076 -214 13140 48
<< metal1 >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18581 3472 18612
rect 1606 18167 3472 18581
rect 3340 18152 3472 18167
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18356 21754 18772
rect 21510 18340 21688 18356
rect 18057 18271 21688 18340
rect 11808 18204 11892 18218
rect 3340 18086 7634 18152
rect 9808 18202 11892 18204
rect 9808 18168 11900 18202
rect 9808 18048 10748 18168
rect 11446 18048 11900 18168
rect 12596 18198 13994 18224
rect 12170 18076 12230 18166
rect 9808 18032 11900 18048
rect 12596 18056 13192 18198
rect 13956 18056 13994 18198
rect 12116 17986 12292 18028
rect 12596 18026 13994 18056
rect 12116 17430 12142 17986
rect 12266 17430 12292 17986
rect 14492 17600 14534 17698
rect 14492 17508 14720 17600
rect 12116 17378 12292 17430
rect 12178 17270 12372 17307
rect 12178 17166 12210 17270
rect 12338 17166 12372 17270
rect 12178 17088 12372 17166
rect 778 16970 23794 17088
rect 778 16960 21572 16970
rect 22312 16960 23794 16970
rect 974 9274 1388 16780
rect 894 9218 1388 9274
rect 892 8944 1388 9218
rect 1582 16688 1986 16710
rect 1582 16576 2556 16688
rect 1582 8950 1692 16576
rect 1838 16496 2556 16576
rect 1838 14602 1986 16496
rect 1838 14368 2640 14602
rect 1838 10470 1986 14368
rect 1838 10236 2708 10470
rect 1838 8950 1986 10236
rect 892 8878 1314 8944
rect 1582 8878 1986 8950
rect 892 8804 1296 8878
rect 892 8592 3720 8804
rect 894 8338 1314 8592
rect 1582 8396 1986 8506
rect 894 696 1006 8338
rect 1214 696 1314 8338
rect 894 584 1314 696
rect 1430 8378 2048 8396
rect 1430 8334 2822 8378
rect 1430 8294 1692 8334
rect 1758 8294 2822 8334
rect 1430 8044 2822 8294
rect 1430 516 2048 8044
rect 2356 6676 2950 6878
rect 12178 684 12372 16960
rect 23220 16664 23636 16916
rect 22720 16330 23090 16482
rect 23220 16424 23736 16664
rect 22720 16190 22818 16330
rect 22852 16190 23090 16330
rect 22720 7934 23090 16190
rect 23266 16412 23736 16424
rect 23266 8756 23332 16412
rect 23638 8756 23736 16412
rect 23266 8582 23736 8756
rect 23538 7956 23636 8582
rect 22614 7888 23090 7934
rect 22614 7792 23004 7888
rect 21734 6674 22524 6954
rect 22614 6286 22698 7792
rect 21712 6004 22698 6286
rect 12182 578 12216 684
rect 12334 578 12368 684
rect 12182 552 12368 578
rect 11996 400 12108 442
rect 3334 182 5004 194
rect 3286 86 5720 182
rect 3286 -36 10302 86
rect 3286 -68 5720 -36
rect 3286 -288 3390 -68
rect 4410 -288 5720 -68
rect 11996 -176 12022 400
rect 12098 -176 12108 400
rect 11996 -196 12108 -176
rect 12358 416 12470 452
rect 12358 -160 12378 416
rect 12454 -160 12470 416
rect 22614 278 22698 6004
rect 22980 278 23004 7792
rect 12358 -186 12470 -160
rect 13016 48 13168 112
rect 22614 110 23004 278
rect 3286 -354 5720 -288
rect 13016 -214 13076 48
rect 13140 -214 13168 48
rect 13016 -312 13168 -214
rect 14208 64 21288 92
rect 14208 -6 20460 64
rect 23202 24 23636 7956
rect 14208 -60 21208 -6
rect 23202 -32 23320 24
rect 14208 -252 19322 -60
rect 21026 -252 21208 -60
rect 12148 -352 12324 -348
rect 12148 -406 12160 -352
rect 12304 -406 12324 -352
rect 12148 -412 12324 -406
rect 13024 -518 13154 -312
rect 14208 -324 21208 -252
rect 19236 -328 21208 -324
rect 23200 -300 23320 -32
rect 23544 -300 23636 24
rect 23200 -386 23636 -300
rect 11518 -539 12126 -518
rect 12306 -539 13334 -518
rect 1278 -669 23744 -539
rect 1640 -912 2170 -868
rect 12976 -910 22452 -896
rect 1640 -948 12234 -912
rect 1640 -980 2170 -948
rect 1640 -2232 1734 -980
rect 2100 -2232 2170 -980
rect 12198 -1468 12234 -948
rect 12976 -928 22780 -910
rect 12976 -932 22422 -928
rect 12546 -1533 12548 -1460
rect 12654 -1486 12690 -1460
rect 12976 -1524 13012 -932
rect 22348 -1916 22422 -932
rect 22738 -1916 22780 -928
rect 22348 -1978 22780 -1916
rect 1640 -2308 2170 -2232
rect 23200 -2330 23636 -910
rect 23210 -4402 23598 -2330
rect 23200 -4756 23636 -4402
rect 13648 -5192 23636 -4756
<< via1 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 10748 18048 11446 18168
rect 13192 18056 13956 18198
rect 12142 17430 12266 17986
rect 3390 -288 4410 -68
rect 12022 -176 12098 400
rect 12378 -160 12454 416
rect 19322 -252 21026 -60
rect 12160 -406 12304 -352
rect 23320 -300 23544 24
rect 1734 -2232 2100 -980
rect 22422 -1916 22738 -928
<< metal2 >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
rect 10708 18168 11484 18202
rect 10708 18048 10748 18168
rect 11446 18048 11484 18168
rect 10708 18020 11484 18048
rect 13150 18198 14006 18228
rect 13150 18056 13192 18198
rect 13956 18056 14006 18198
rect 13150 18030 14006 18056
rect 12114 17986 12298 18028
rect 12114 17510 12142 17986
rect 12108 17430 12142 17510
rect 12266 17430 12298 17986
rect 12108 17380 12298 17430
rect 12108 17100 12288 17380
rect 778 17036 23284 17100
rect 10266 15868 14172 15920
rect 10308 13784 14220 13836
rect 10336 11702 14134 11754
rect 10426 9616 14124 9668
rect 10388 7530 14150 7582
rect 10400 5448 14162 5500
rect 10362 3360 14262 3412
rect 10436 1276 14166 1328
rect 11996 400 12108 442
rect 3286 -68 4540 -24
rect 3286 -288 3390 -68
rect 4410 -288 4540 -68
rect 11996 -176 12022 400
rect 12098 -176 12108 400
rect 11996 -196 12108 -176
rect 12358 416 12470 452
rect 12358 -160 12378 416
rect 12454 -160 12470 416
rect 23208 24 23634 80
rect 12358 -186 12470 -160
rect 19270 -60 21100 -16
rect 3286 -290 3392 -288
rect 4404 -290 4540 -288
rect 3286 -354 4540 -290
rect 19270 -252 19322 -60
rect 21026 -252 21100 -60
rect 19270 -326 21100 -252
rect 23208 -300 23320 24
rect 23544 -300 23634 24
rect 12148 -352 12324 -348
rect 12148 -406 12160 -352
rect 12304 -406 12324 -352
rect 23208 -370 23634 -300
rect 12148 -412 12324 -406
rect 12172 -526 12278 -412
rect 796 -766 23680 -526
rect 1640 -980 2170 -868
rect 1640 -2232 1734 -980
rect 2100 -2232 2170 -980
rect 22348 -928 22780 -872
rect 22348 -1916 22422 -928
rect 22738 -1916 22780 -928
rect 22348 -1978 22780 -1916
rect 1640 -2308 2170 -2232
<< via2 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 10748 18048 11446 18168
rect 13192 18056 13956 18198
rect 3390 -288 4410 -68
rect 12022 -176 12098 400
rect 12378 -160 12454 416
rect 3392 -290 4404 -288
rect 19322 -252 21026 -60
rect 23320 -300 23544 24
rect 1734 -2232 2100 -980
rect 22422 -1916 22738 -928
<< metal3 >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
rect 10708 18168 11484 18202
rect 10708 18048 10748 18168
rect 11446 18048 11484 18168
rect 10708 18020 11484 18048
rect 13150 18198 14006 18228
rect 13150 18056 13192 18198
rect 13956 18056 14006 18198
rect 13150 18030 14006 18056
rect 1646 17280 10212 17800
rect 1646 -868 2166 17280
rect 11796 15580 11968 17674
rect 12444 15570 12616 17664
rect 15074 17546 22766 17966
rect 11996 400 12108 442
rect 11996 124 12022 400
rect 8604 112 12022 124
rect 8592 68 12022 112
rect 3286 -68 4540 -24
rect 3286 -288 3390 -68
rect 4410 -288 4540 -68
rect 8592 -154 8658 68
rect 10706 -154 12022 68
rect 8592 -176 12022 -154
rect 12098 -176 12108 400
rect 8592 -184 12108 -176
rect 8592 -196 10830 -184
rect 11996 -196 12108 -184
rect 12358 416 12470 452
rect 12358 -160 12378 416
rect 12454 118 12470 416
rect 14010 118 17022 130
rect 12454 68 17022 118
rect 12454 -128 14114 68
rect 16924 -128 17022 68
rect 12454 -160 17022 -128
rect 12358 -178 17022 -160
rect 19270 -60 21100 -16
rect 12358 -186 12470 -178
rect 3286 -290 3392 -288
rect 4404 -290 4540 -288
rect 3286 -354 4540 -290
rect 19270 -252 19322 -60
rect 21026 -252 21100 -60
rect 19270 -326 21100 -252
rect 1640 -980 2170 -868
rect 1640 -2232 1734 -980
rect 2100 -1816 2170 -980
rect 22346 -872 22766 17546
rect 23208 24 23634 80
rect 23208 -300 23320 24
rect 23544 -300 23634 24
rect 23208 -370 23634 -300
rect 22346 -928 22780 -872
rect 15760 -1694 15828 -1580
rect 2100 -2232 8918 -1816
rect 22346 -1916 22422 -928
rect 22738 -1916 22780 -928
rect 22346 -1956 22780 -1916
rect 1640 -2308 8918 -2232
rect 1646 -2336 8918 -2308
rect 16944 -1978 22780 -1956
rect 16944 -2330 22766 -1978
rect 16944 -2376 22016 -2330
rect 12520 -7844 12606 -7576
<< via3 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 10748 18048 11446 18168
rect 13192 18056 13956 18198
rect 3390 -288 4410 -68
rect 8658 -154 10706 68
rect 14114 -128 16924 68
rect 3392 -290 4404 -288
rect 19322 -252 21026 -60
rect 23320 -300 23544 24
<< metal4 >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 12596 18198 14680 18216
rect 3340 18086 7634 18152
rect 9804 18168 11832 18190
rect 9804 18048 10748 18168
rect 11446 18048 11832 18168
rect 9804 18018 11832 18048
rect 12596 18056 13192 18198
rect 13956 18056 14680 18198
rect 12596 18026 14680 18056
rect 1358 -4701 2016 1587
rect 16482 130 17004 133
rect 8604 112 9236 126
rect 8592 68 10830 112
rect 3286 -68 4540 -24
rect 3286 -288 3390 -68
rect 4410 -288 4540 -68
rect 8592 -154 8658 68
rect 10706 -154 10830 68
rect 8592 -196 10830 -154
rect 14010 68 17022 130
rect 14010 -128 14114 68
rect 16924 -128 17022 68
rect 19270 -26 21100 -16
rect 22504 -26 23162 1763
rect 14010 -178 17022 -128
rect 19236 -60 23162 -26
rect 3286 -290 3392 -288
rect 4404 -290 4540 -288
rect 3286 -354 4540 -290
rect 3288 -4701 4518 -354
rect 8604 -2440 9236 -196
rect 16482 -1856 17004 -178
rect 19236 -252 19322 -60
rect 21026 -252 23162 -60
rect 19236 -294 23162 -252
rect 19270 -326 21100 -294
rect 22504 -386 23162 -294
rect 23256 24 23628 76
rect 23256 -300 23320 24
rect 23560 -300 23628 24
rect 23256 -370 23628 -300
rect 22504 -596 22868 -386
rect 22504 -750 22922 -596
rect 22504 -2330 23162 -750
rect 1358 -5352 11601 -4701
rect 1358 -5359 7050 -5352
rect 11190 -5359 11601 -5352
rect 11190 -5624 11584 -5359
<< via4 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 23320 -300 23544 24
rect 23544 -300 23560 24
<< metal5 >>
rect 20959 18861 23756 18883
rect 18057 18772 23756 18861
rect 764 18650 3585 18679
rect 764 18612 7634 18650
rect 764 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 23756 18772
rect 18057 18271 23756 18340
rect 20743 18203 23756 18271
rect 764 18086 7634 18152
rect 764 18035 4377 18086
rect 764 18021 3585 18035
rect 764 17960 1422 18021
rect 778 16744 1422 17960
rect 764 14595 1422 16744
rect 23098 14615 23756 18203
rect 23043 24 23633 1129
rect 23043 -300 23320 24
rect 23560 -300 23633 24
rect 23043 -4695 23633 -300
rect 13677 -5285 23633 -4695
use capacitors_5  capacitors_5_0
timestamp 1699177610
transform 1 0 2736 0 1 14838
box -1972 -14958 10096 2068
use capacitors_5  capacitors_5_1
timestamp 1699177610
transform -1 0 21784 0 1 14844
box -1972 -14958 10096 2068
use clock  clock_0
timestamp 1699103691
transform 0 -1 12414 1 0 -7452
box -410 -1832 6030 1274
use nmos_diode2  nmos_diode2_0
timestamp 1699103691
transform 1 0 11416 0 1 576
box -46 -1200 1896 182
use nmos_dnw3  nmos_dnw3_0
timestamp 1699103691
transform 1 0 11936 0 1 16204
box -424 892 1176 2258
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_0
timestamp 1699103691
transform -1 0 16844 0 1 -2266
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_1
timestamp 1699103691
transform 1 0 8830 0 1 -2176
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_4
timestamp 1699103691
transform -1 0 9516 0 1 18074
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_5
timestamp 1699103691
transform 1 0 15220 0 1 18046
box -1086 -940 1086 940
use sky130_fd_pr__nfet_01v8_NJGC8F  sky130_fd_pr__nfet_01v8_NJGC8F_0
timestamp 1699103691
transform 0 1 1358 -1 0 12825
box -3869 -130 3869 130
use sky130_fd_pr__nfet_01v8_NJGC8F  sky130_fd_pr__nfet_01v8_NJGC8F_1
timestamp 1699103691
transform 0 1 23234 -1 0 4047
box -3869 -130 3869 130
use sky130_fd_pr__pfet_01v8_4RPJ49  sky130_fd_pr__pfet_01v8_4RPJ49_0
timestamp 1699103691
transform 0 -1 1472 1 0 4485
box -3905 -142 3905 142
use sky130_fd_pr__pfet_01v8_4RPJ49  sky130_fd_pr__pfet_01v8_4RPJ49_1
timestamp 1699103691
transform 0 1 23042 -1 0 12489
box -3905 -142 3905 142
<< labels >>
rlabel metal1 12198 18156 12198 18156 1 vin
port 3 n
rlabel metal1 12266 16974 12266 16974 1 vs
port 4 n
rlabel space 11822 15478 11822 15478 1 input1
port 5 n
rlabel space 12698 15690 12698 15690 1 input2
port 6 n
rlabel metal2 12044 15902 12044 15902 1 in1
port 7 n
rlabel metal2 12868 13820 12868 13820 1 in2
port 8 n
rlabel metal2 12816 11730 12816 11730 1 in3
port 9 n
rlabel metal2 12818 9640 12818 9640 1 in4
port 10 n
rlabel metal2 12646 7556 12646 7556 1 in5
port 11 n
rlabel metal2 12808 5478 12808 5478 1 in6
port 12 n
rlabel metal2 12078 3396 12078 3396 1 in7
port 13 n
rlabel metal2 12050 1306 12050 1306 1 in8
port 14 n
rlabel metal3 10706 -184 12022 124 1 input1
port 15 n
rlabel metal3 13376 -92 13376 -92 1 input2
port 16 n
rlabel metal2 12228 -446 12228 -446 1 out
port 17 n
rlabel metal1 11410 -936 11410 -936 1 clk
port 18 n
rlabel metal1 13184 -910 13184 -910 1 clkb
port 19 n
rlabel metal3 12564 -7798 12564 -7798 1 clk_in
port 20 n
rlabel metal4 10632 18112 10632 18112 1 g1
port 21 n
rlabel metal4 14056 18118 14056 18118 1 g2
port 22 n
<< end >>
