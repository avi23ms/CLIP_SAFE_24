magic
tech sky130A
magscale 1 2
timestamp 1699103691
<< nmos >>
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
<< ndiff >>
rect -413 30 -351 42
rect -413 -30 -401 30
rect -367 -30 -351 30
rect -413 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 413 42
rect 351 -30 367 30
rect 401 -30 413 30
rect 351 -42 413 -30
<< ndiffc >>
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
<< poly >>
rect -273 114 -207 130
rect -273 80 -257 114
rect -223 80 -207 114
rect -351 42 -321 68
rect -273 64 -207 80
rect -81 114 -15 130
rect -81 80 -65 114
rect -31 80 -15 114
rect -255 42 -225 64
rect -159 42 -129 68
rect -81 64 -15 80
rect 111 114 177 130
rect 111 80 127 114
rect 161 80 177 114
rect -63 42 -33 64
rect 33 42 63 68
rect 111 64 177 80
rect 303 114 369 130
rect 303 80 319 114
rect 353 80 369 114
rect 129 42 159 64
rect 225 42 255 68
rect 303 64 369 80
rect 321 42 351 64
rect -351 -64 -321 -42
rect -369 -80 -303 -64
rect -255 -68 -225 -42
rect -159 -64 -129 -42
rect -369 -114 -353 -80
rect -319 -114 -303 -80
rect -369 -130 -303 -114
rect -177 -80 -111 -64
rect -63 -68 -33 -42
rect 33 -64 63 -42
rect -177 -114 -161 -80
rect -127 -114 -111 -80
rect -177 -130 -111 -114
rect 15 -80 81 -64
rect 129 -68 159 -42
rect 225 -64 255 -42
rect 15 -114 31 -80
rect 65 -114 81 -80
rect 15 -130 81 -114
rect 207 -80 273 -64
rect 321 -68 351 -42
rect 207 -114 223 -80
rect 257 -114 273 -80
rect 207 -130 273 -114
<< polycont >>
rect -257 80 -223 114
rect -65 80 -31 114
rect 127 80 161 114
rect 319 80 353 114
rect -353 -114 -319 -80
rect -161 -114 -127 -80
rect 31 -114 65 -80
rect 223 -114 257 -80
<< locali >>
rect -273 80 -257 114
rect -223 80 -207 114
rect -81 80 -65 114
rect -31 80 -15 114
rect 111 80 127 114
rect 161 80 177 114
rect 303 80 319 114
rect 353 80 369 114
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect -369 -114 -353 -80
rect -319 -114 -303 -80
rect -177 -114 -161 -80
rect -127 -114 -111 -80
rect 15 -114 31 -80
rect 65 -114 81 -80
rect 207 -114 223 -80
rect 257 -114 273 -80
<< viali >>
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
<< metal1 >>
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
