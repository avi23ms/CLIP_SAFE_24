magic
tech sky130A
magscale 1 2
timestamp 1698902756
<< pwell >>
rect 554 1146 591 1291
rect 1630 1192 1660 1286
rect 1958 1044 2056 1226
rect 3476 932 3550 1002
rect 4364 918 4550 1024
rect 4364 866 4742 918
rect 4542 850 4742 866
<< poly >>
rect 234 2243 264 2244
rect 234 2213 357 2243
rect 234 2184 264 2213
rect 2944 2053 2974 2122
rect 2845 2023 2974 2053
rect 3898 1084 3955 1114
rect 3925 1011 3955 1084
<< locali >>
rect 4644 2372 4684 2374
rect 223 2340 4950 2372
rect 223 2337 3600 2340
rect 4928 2296 4950 2340
rect 3627 2295 4950 2296
rect 223 2235 4950 2295
rect 1279 2106 1347 2235
rect 2435 2098 2503 2235
rect 3448 2228 4950 2235
rect 4644 1870 4684 2228
rect 1101 1688 1524 1725
rect 2262 1689 2685 1726
rect 1132 1172 1549 1215
rect 2287 1199 2706 1208
rect 2287 1166 2707 1199
rect 1301 998 1376 1096
rect 2464 998 2532 1100
rect 226 986 3476 998
rect 226 932 3558 986
rect 3790 914 3888 974
rect 4542 914 4742 918
rect 3558 909 4742 914
rect 3558 890 4179 909
rect 215 869 4179 890
rect 4541 869 4742 909
rect 215 850 4742 869
rect 3802 848 3890 850
<< viali >>
rect 3600 2337 4928 2340
rect 218 2296 4928 2337
rect 218 2295 3627 2296
rect 215 890 3558 932
rect 4179 869 4541 909
<< metal1 >>
rect -25 2343 305 2349
rect 3482 2343 4950 2372
rect -25 2340 4950 2343
rect -25 2337 3600 2340
rect -25 2307 218 2337
rect -25 1195 17 2307
rect 160 2299 218 2307
rect 206 2295 218 2299
rect 4928 2296 4950 2340
rect 3627 2295 4950 2296
rect 206 2234 4950 2295
rect 206 2232 2156 2234
rect 2218 2232 4950 2234
rect 206 2228 248 2232
rect 1589 2230 1621 2232
rect 3482 2228 4950 2232
rect 3562 2224 3602 2228
rect 124 2126 984 2174
rect 124 2100 214 2126
rect 2795 2107 3623 2157
rect 124 1738 172 2100
rect 222 2014 852 2064
rect 2832 2008 3474 2060
rect 1556 1754 1638 1767
rect 328 1738 338 1742
rect 124 1690 338 1738
rect 328 1675 338 1690
rect 393 1675 403 1742
rect 514 1716 591 1753
rect 514 1708 551 1716
rect 552 1708 591 1716
rect 514 1671 591 1708
rect 552 1636 591 1671
rect 714 1668 724 1735
rect 779 1668 789 1735
rect 898 1666 976 1753
rect 1556 1681 1571 1754
rect 1639 1681 1649 1754
rect 1556 1667 1638 1681
rect 451 1279 480 1632
rect 554 1441 591 1636
rect 814 1580 824 1632
rect 886 1580 896 1632
rect 943 1442 976 1666
rect 1679 1442 1712 1850
rect 1759 1665 1842 1702
rect 1805 1636 1842 1665
rect 1806 1629 1842 1636
rect 1806 1576 1844 1629
rect 1806 1572 1842 1576
rect 943 1441 1712 1442
rect 552 1411 1712 1441
rect 354 1195 364 1203
rect -25 1153 364 1195
rect 354 1136 364 1153
rect 419 1136 429 1203
rect 554 1146 591 1411
rect 943 1409 1712 1411
rect 825 1269 835 1321
rect 897 1269 907 1321
rect 746 1133 756 1200
rect 811 1133 821 1200
rect 943 1145 976 1409
rect 1600 1194 1668 1242
rect 1805 1226 1842 1572
rect 1600 1134 1674 1194
rect 1726 1146 1842 1226
rect 1973 1241 2007 1762
rect 2078 1442 2111 1844
rect 2140 1673 2150 1761
rect 2218 1673 2228 1761
rect 2835 1759 2868 1770
rect 2835 1659 2876 1759
rect 2999 1665 3009 1732
rect 3064 1665 3074 1732
rect 2835 1442 2868 1659
rect 2906 1576 2916 1628
rect 2981 1576 2991 1628
rect 2078 1440 2868 1442
rect 3210 1440 3247 1761
rect 3387 1673 3397 1740
rect 3452 1722 3462 1740
rect 3573 1722 3623 2107
rect 3452 1673 3624 1722
rect 3392 1672 3624 1673
rect 2078 1410 3247 1440
rect 2078 1409 2868 1410
rect 1973 1219 2046 1241
rect 2835 1240 2868 1409
rect 2934 1268 2944 1320
rect 3009 1268 3019 1320
rect -95 1061 507 1100
rect 280 956 290 997
rect 223 940 290 956
rect 361 956 371 997
rect 1608 956 1636 1134
rect 1726 1100 1822 1146
rect 1954 1140 1964 1219
rect 2037 1140 2047 1219
rect 2194 1199 2230 1238
rect 2188 1139 2239 1199
rect 2835 1143 2910 1240
rect 3210 1239 3247 1410
rect 3330 1273 3370 1621
rect 3031 1147 3041 1214
rect 3096 1147 3106 1214
rect 1726 1062 2066 1100
rect 1768 1054 2066 1062
rect 2194 956 2230 1139
rect 3210 1128 3290 1239
rect 3416 1147 3426 1214
rect 3481 1195 3491 1214
rect 3481 1193 3521 1195
rect 3654 1194 3694 2228
rect 3923 1749 4027 1763
rect 3923 1564 3937 1749
rect 4015 1564 4027 1749
rect 4157 1568 4197 2228
rect 3923 1554 4027 1564
rect 4340 1559 4419 1765
rect 4546 1569 4586 2228
rect 4348 1514 4391 1559
rect 4348 1510 4511 1514
rect 4045 1475 4511 1510
rect 4348 1470 4511 1475
rect 3654 1193 3752 1194
rect 3481 1154 3752 1193
rect 3481 1153 3620 1154
rect 3481 1147 3491 1153
rect 3332 1096 3666 1101
rect 2970 1064 3666 1096
rect 3712 1074 3752 1154
rect 2970 1058 3403 1064
rect 3474 986 3615 999
rect 3474 956 3484 986
rect 361 940 3484 956
rect 223 938 3484 940
rect 203 932 3484 938
rect 3541 956 3615 986
rect 3802 974 3878 1258
rect 3541 932 3573 956
rect 203 890 215 932
rect 3558 912 3573 932
rect 3790 914 3888 974
rect 3920 972 3960 1222
rect 4348 1148 4391 1470
rect 4096 1062 4965 1103
rect 4614 1059 4965 1062
rect 4366 1024 4545 1025
rect 4364 920 4550 1024
rect 4276 918 4550 920
rect 4276 915 4742 918
rect 3790 912 3892 914
rect 4167 912 4742 915
rect 3558 909 4742 912
rect 3558 890 4179 909
rect 203 884 4179 890
rect 223 869 4179 884
rect 4541 869 4742 909
rect 223 853 4742 869
rect 3412 850 4742 853
rect 3412 848 4677 850
<< via1 >>
rect 338 1675 393 1742
rect 724 1668 779 1735
rect 1571 1681 1639 1754
rect 824 1580 886 1632
rect 364 1136 419 1203
rect 835 1269 897 1321
rect 756 1133 811 1200
rect 2150 1673 2218 1761
rect 3009 1665 3064 1732
rect 2916 1576 2981 1628
rect 3397 1673 3452 1740
rect 2944 1268 3009 1320
rect 290 940 361 997
rect 1964 1140 2037 1219
rect 3041 1147 3096 1214
rect 3426 1147 3481 1214
rect 3937 1564 4015 1749
rect 3484 932 3541 986
<< metal2 >>
rect 1551 2333 2187 2337
rect 3736 2333 4011 2344
rect 1551 2307 4011 2333
rect 1551 2304 3921 2307
rect 1551 2296 3868 2304
rect 829 1855 859 1860
rect -125 1845 869 1855
rect -125 1814 875 1845
rect -125 1813 869 1814
rect 338 1742 393 1752
rect 295 1739 338 1740
rect 216 1696 338 1739
rect 216 992 259 1696
rect 295 1695 338 1696
rect 319 1691 338 1695
rect 724 1735 779 1745
rect 393 1691 724 1727
rect 338 1665 393 1675
rect 724 1658 779 1668
rect 829 1642 859 1813
rect 1551 1767 1588 2296
rect 2150 1771 2187 2296
rect 1551 1764 1638 1767
rect 1551 1754 1639 1764
rect 1551 1681 1571 1754
rect 1551 1671 1639 1681
rect 2150 1761 2218 1771
rect 3974 1763 4011 2307
rect 1551 1667 1638 1671
rect 2150 1663 2218 1673
rect 3009 1732 3064 1742
rect 3397 1740 3452 1750
rect 3064 1682 3397 1718
rect 3009 1655 3064 1665
rect 3923 1749 4027 1763
rect 3452 1676 3618 1718
rect 3397 1663 3452 1673
rect 824 1632 886 1642
rect 824 1570 886 1580
rect 2916 1630 2981 1638
rect 2916 1628 2982 1630
rect 2981 1576 2982 1628
rect 832 1331 867 1570
rect 2916 1566 2982 1576
rect 832 1321 897 1331
rect 2946 1330 2982 1566
rect 832 1278 835 1321
rect 835 1259 897 1269
rect 2944 1320 3009 1330
rect 2944 1258 3009 1268
rect 1964 1226 2037 1229
rect 1958 1219 2056 1226
rect 364 1203 419 1213
rect 349 1143 364 1179
rect 756 1200 811 1210
rect 419 1143 756 1179
rect 364 1126 419 1136
rect 756 1123 811 1133
rect 1958 1140 1964 1219
rect 2037 1140 2056 1219
rect 3041 1214 3096 1224
rect 3036 1157 3041 1193
rect 1958 1044 2056 1140
rect 3426 1214 3481 1224
rect 3096 1157 3426 1193
rect 3041 1137 3096 1147
rect 3481 1157 3487 1193
rect 3426 1137 3481 1147
rect 306 1007 349 1014
rect 290 997 361 1007
rect 216 949 290 992
rect 361 949 363 992
rect 290 930 361 940
rect 1960 858 2056 1044
rect 3576 1029 3618 1676
rect 3923 1564 3937 1749
rect 4015 1564 4027 1749
rect 3923 1554 4027 1564
rect 3477 1002 3618 1029
rect 3476 986 3618 1002
rect 3476 932 3484 986
rect 3541 939 3618 986
rect 3541 932 3550 939
rect 3484 922 3541 932
rect -158 762 2056 858
<< via2 >>
rect 1964 1140 2037 1219
<< metal3 >>
rect 1948 1219 2048 1230
rect 1948 1140 1964 1219
rect 2037 1140 2048 1219
rect 1948 1134 2048 1140
use sky130_fd_pr__nfet_01v8_3374R3  sky130_fd_pr__nfet_01v8_3374R3_0
timestamp 1698871184
transform 0 1 4382 1 0 1088
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_GWAZJ9  sky130_fd_pr__nfet_01v8_GWAZJ9_0
timestamp 1698873245
transform 1 0 3199 0 1 2132
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_0
timestamp 1698873245
transform 1 0 585 0 1 2142
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_J7MSU8  sky130_fd_pr__nfet_01v8_J7MSU8_0
timestamp 1698873245
transform 0 -1 3842 1 0 1099
box -173 -130 173 130
use sky130_fd_pr__pfet_01v8_BH9SS5  sky130_fd_pr__pfet_01v8_BH9SS5_0
timestamp 1698787694
transform -1 0 4082 0 -1 1659
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_BH9SS5  sky130_fd_pr__pfet_01v8_BH9SS5_1
timestamp 1698787694
transform 1 0 4468 0 1 1659
box -246 -319 246 319
use sky130_fd_pr__nfet_01v8_SMGLWN  XM1
timestamp 1698155087
transform 1 0 1340 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM2
timestamp 1698155087
transform 1 0 2498 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_PDYTS5  XM3
timestamp 1698869571
transform 1 0 1313 0 1 1866
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_TM5SY6  XM4
timestamp 1698155087
transform 1 0 453 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_PDYTS5  XM5
timestamp 1698869571
transform 1 0 1699 0 1 1866
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_PDYTS5  XM6
timestamp 1698869571
transform 1 0 2085 0 1 1866
box -246 -419 246 419
use sky130_fd_pr__nfet_01v8_SMGLWN  XM7
timestamp 1698155087
transform 1 0 1726 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM8
timestamp 1698155087
transform 1 0 2112 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM10
timestamp 1698155087
transform 1 0 480 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM11
timestamp 1698155087
transform 1 0 866 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_TM5SY6  XM12
timestamp 1698155087
transform 1 0 839 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__nfet_01v8_SMGLWN  XM13
timestamp 1698155087
transform 1 0 2972 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM14
timestamp 1698155087
transform 1 0 3358 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_TM5SY6  XM15
timestamp 1698155087
transform 1 0 2945 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  XM16
timestamp 1698155087
transform 1 0 3331 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_PDYTS5  XM18
timestamp 1698869571
transform 1 0 2471 0 1 1866
box -246 -419 246 419
<< labels >>
rlabel metal1 1405 853 1405 853 5 gnd
rlabel locali 1990 2372 1990 2372 1 Vdd
rlabel metal1 -31 1076 -31 1076 1 vin
rlabel metal2 -68 1827 -68 1827 1 vin2
rlabel metal1 2893 1440 2893 1440 1 Vcm
rlabel metal1 4841 1074 4841 1074 1 Vbias
rlabel metal2 -110 808 -110 808 1 Vb
rlabel metal1 4860 2268 4860 2268 1 Vdd
rlabel metal1 4692 870 4692 870 1 gnd
rlabel metal1 3634 1076 3634 1076 1 Vref
<< end >>
