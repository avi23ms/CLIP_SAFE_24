magic
tech sky130A
magscale 1 2
timestamp 1698205020
<< dnwell >>
rect -254 2142 1076 2232
rect -254 2048 1214 2142
rect -400 2034 1214 2048
rect -418 1130 1302 2034
rect -254 1020 1214 1130
rect -254 906 1076 1020
<< nwell >>
rect -424 2040 1302 2256
rect -424 1130 -252 2040
rect 1072 1132 1302 2040
rect 748 1130 1302 1132
rect -424 896 1302 1130
rect -194 894 1254 896
<< nmos >>
rect 80 1858 110 1942
rect 668 1858 698 1942
rect 0 1200 200 1800
rect 590 1200 790 1800
<< ndiff >>
rect 20 1920 80 1942
rect 20 1882 30 1920
rect 64 1882 80 1920
rect 20 1858 80 1882
rect 110 1928 172 1942
rect 110 1872 124 1928
rect 158 1872 172 1928
rect 110 1858 172 1872
rect 606 1928 668 1942
rect 606 1872 620 1928
rect 654 1872 668 1928
rect 606 1858 668 1872
rect 698 1920 758 1942
rect 698 1882 714 1920
rect 748 1882 758 1920
rect 698 1858 758 1882
rect -110 1770 0 1800
rect -110 1230 -90 1770
rect -40 1230 0 1770
rect -110 1200 0 1230
rect 200 1770 310 1800
rect 200 1230 230 1770
rect 280 1230 310 1770
rect 200 1200 310 1230
rect 480 1770 590 1800
rect 480 1230 510 1770
rect 560 1230 590 1770
rect 480 1200 590 1230
rect 790 1770 900 1800
rect 790 1230 830 1770
rect 880 1230 900 1770
rect 790 1200 900 1230
<< ndiffc >>
rect 30 1882 64 1920
rect 124 1872 158 1928
rect 620 1872 654 1928
rect 714 1882 748 1920
rect -90 1230 -40 1770
rect 230 1230 280 1770
rect 510 1230 560 1770
rect 830 1230 880 1770
<< psubdiff >>
rect -66 1920 20 1942
rect -66 1882 -40 1920
rect -6 1882 20 1920
rect -66 1858 20 1882
rect 758 1920 844 1942
rect 758 1882 784 1920
rect 818 1882 844 1920
rect 758 1858 844 1882
rect -220 1770 -110 1800
rect -220 1230 -190 1770
rect -140 1230 -110 1770
rect -220 1200 -110 1230
rect 900 1770 1010 1800
rect 900 1230 930 1770
rect 980 1230 1010 1770
rect 900 1200 1010 1230
<< nsubdiff >>
rect 912 2216 1004 2220
rect -210 2190 -122 2210
rect 910 2200 1004 2216
rect -210 2108 -184 2190
rect -146 2108 -122 2190
rect 908 2196 1004 2200
rect 908 2112 932 2196
rect -210 2078 -122 2108
rect 910 2102 932 2112
rect 980 2102 1004 2196
rect 910 2078 1004 2102
<< psubdiffcont >>
rect -40 1882 -6 1920
rect 784 1882 818 1920
rect -190 1230 -140 1770
rect 930 1230 980 1770
<< nsubdiffcont >>
rect -184 2108 -146 2190
rect 932 2102 980 2196
<< poly >>
rect 80 1942 110 1972
rect 668 1942 698 1972
rect 80 1826 110 1858
rect 668 1826 698 1858
rect 0 1800 200 1826
rect 590 1800 790 1826
rect 0 1172 200 1200
rect 590 1174 790 1200
<< locali >>
rect 912 2216 1004 2220
rect -210 2190 -122 2210
rect 910 2200 1004 2216
rect -210 2108 -184 2190
rect -146 2108 -122 2190
rect 908 2196 1004 2200
rect 908 2112 932 2196
rect -210 2070 -122 2108
rect 910 2102 932 2112
rect 980 2102 1004 2196
rect 910 2078 1004 2102
rect -42 1924 74 1936
rect -42 1878 -40 1924
rect 64 1878 74 1924
rect -42 1864 74 1878
rect 114 1934 170 1944
rect 114 1866 124 1934
rect 158 1866 170 1934
rect 114 1854 170 1866
rect 608 1934 664 1944
rect 608 1866 620 1934
rect 654 1866 664 1934
rect 608 1854 664 1866
rect 704 1924 820 1936
rect 704 1878 714 1924
rect 818 1878 820 1924
rect 704 1864 820 1878
rect -122 1790 -2 1804
rect -210 1770 -2 1790
rect -210 1230 -190 1770
rect -140 1230 -90 1770
rect -40 1230 -2 1770
rect 202 1770 302 1796
rect 202 1768 230 1770
rect 202 1734 228 1768
rect -210 1210 -2 1230
rect 210 1234 228 1734
rect 280 1734 302 1770
rect 480 1790 578 1800
rect 790 1790 910 1818
rect 480 1770 580 1790
rect 480 1766 510 1770
rect 480 1758 508 1766
rect 210 1230 230 1234
rect 280 1230 300 1734
rect 210 1210 300 1230
rect 490 1234 508 1758
rect 490 1230 510 1234
rect 560 1230 580 1770
rect 490 1210 580 1230
rect 790 1770 1000 1790
rect 790 1230 830 1770
rect 880 1230 930 1770
rect 980 1230 1000 1770
rect 790 1210 1000 1230
rect -122 1190 -2 1210
rect 790 1204 910 1210
<< viali >>
rect -184 2108 -146 2190
rect 932 2102 980 2196
rect -40 1920 64 1924
rect -40 1882 -6 1920
rect -6 1882 30 1920
rect 30 1882 64 1920
rect -40 1878 64 1882
rect 124 1928 158 1934
rect 124 1872 158 1928
rect 124 1866 158 1872
rect 620 1928 654 1934
rect 620 1872 654 1928
rect 620 1866 654 1872
rect 714 1920 818 1924
rect 714 1882 748 1920
rect 748 1882 784 1920
rect 784 1882 818 1920
rect 714 1878 818 1882
rect -190 1230 -140 1770
rect 228 1234 230 1768
rect 230 1234 280 1768
rect 508 1234 510 1766
rect 510 1234 560 1766
rect 930 1230 980 1770
<< metal1 >>
rect -208 2324 1004 2410
rect -208 2322 20 2324
rect 96 2322 704 2324
rect 780 2322 1004 2324
rect -208 2210 -120 2322
rect 916 2216 1004 2322
rect -210 2190 -120 2210
rect -210 2108 -184 2190
rect -146 2152 -120 2190
rect 910 2196 1004 2216
rect -146 2108 -122 2152
rect -210 2094 -122 2108
rect 910 2102 932 2196
rect 980 2120 1004 2196
rect 980 2102 1000 2120
rect -210 2052 -126 2094
rect 910 2084 1000 2102
rect 908 2056 1000 2084
rect -210 1930 -122 2052
rect -36 1930 74 1936
rect -210 1924 74 1930
rect -210 1878 -40 1924
rect 64 1878 74 1924
rect -210 1868 74 1878
rect -210 1802 -122 1868
rect -36 1864 74 1868
rect 112 1934 170 1946
rect 112 1866 124 1934
rect 158 1866 170 1934
rect 112 1854 170 1866
rect 608 1934 666 1946
rect 608 1866 620 1934
rect 654 1866 666 1934
rect 608 1854 666 1866
rect 704 1930 814 1936
rect 910 1930 1000 2056
rect 704 1924 1000 1930
rect 704 1878 714 1924
rect 818 1878 1000 1924
rect 704 1868 1000 1878
rect 704 1864 814 1868
rect -210 1770 -120 1802
rect -210 1230 -190 1770
rect -140 1230 -120 1770
rect -210 1190 -120 1230
rect 200 1772 312 1802
rect 200 1230 210 1772
rect 302 1230 312 1772
rect 480 1772 590 1800
rect 480 1269 494 1772
rect 200 1202 312 1230
rect 479 1230 494 1269
rect 576 1230 590 1772
rect 910 1770 1000 1868
rect 910 1380 930 1770
rect 479 1202 590 1230
rect 908 1230 930 1380
rect 980 1230 1000 1770
rect 908 1220 1000 1230
rect 210 1190 300 1202
rect 479 1190 569 1202
rect 908 1190 998 1220
<< via1 >>
rect 210 1768 302 1772
rect 210 1234 228 1768
rect 228 1234 280 1768
rect 280 1234 302 1768
rect 210 1230 302 1234
rect 494 1766 576 1772
rect 494 1234 508 1766
rect 508 1234 560 1766
rect 560 1234 576 1766
rect 494 1230 576 1234
<< metal2 >>
rect 200 1772 312 1802
rect 200 1230 210 1772
rect 302 1230 312 1772
rect 200 1202 312 1230
rect 480 1772 590 1800
rect 480 1230 494 1772
rect 576 1230 590 1772
rect 480 1202 590 1230
<< via2 >>
rect 210 1230 302 1772
rect 494 1230 576 1772
<< metal3 >>
rect 200 1772 312 1802
rect 200 1230 210 1772
rect 302 1230 312 1772
rect 200 818 312 1230
rect 480 1772 590 1800
rect 480 1230 494 1772
rect 576 1268 590 1772
rect 576 1230 592 1268
rect 480 832 592 1230
<< end >>
