magic
tech sky130A
magscale 1 2
timestamp 1698662012
<< nwell >>
rect 21388 -666 21824 -290
rect 23830 -640 24266 -264
rect 66988 -666 67424 -290
rect 69430 -640 69866 -264
rect 89788 -666 90224 -290
rect 92230 -640 92666 -264
<< nmos >>
rect 21482 -818 21512 -734
rect 21700 -818 21730 -734
rect 23924 -792 23954 -708
rect 24142 -792 24172 -708
rect 67082 -818 67112 -734
rect 67300 -818 67330 -734
rect 69524 -792 69554 -708
rect 69742 -792 69772 -708
rect 89882 -818 89912 -734
rect 90100 -818 90130 -734
rect 92324 -792 92354 -708
rect 92542 -792 92572 -708
<< pmos >>
rect 21482 -604 21512 -352
rect 21700 -604 21730 -352
rect 23924 -578 23954 -326
rect 24142 -578 24172 -326
rect 67082 -604 67112 -352
rect 67300 -604 67330 -352
rect 69524 -578 69554 -326
rect 69742 -578 69772 -326
rect 89882 -604 89912 -352
rect 90100 -604 90130 -352
rect 92324 -578 92354 -326
rect 92542 -578 92572 -326
<< ndiff >>
rect 23866 -720 23924 -708
rect 21424 -746 21482 -734
rect 21424 -806 21436 -746
rect 21470 -806 21482 -746
rect 21424 -818 21482 -806
rect 21512 -746 21570 -734
rect 21512 -806 21524 -746
rect 21558 -806 21570 -746
rect 21512 -818 21570 -806
rect 21642 -746 21700 -734
rect 21642 -806 21654 -746
rect 21688 -806 21700 -746
rect 21642 -818 21700 -806
rect 21730 -746 21788 -734
rect 21730 -806 21742 -746
rect 21776 -806 21788 -746
rect 23866 -780 23878 -720
rect 23912 -780 23924 -720
rect 23866 -792 23924 -780
rect 23954 -720 24012 -708
rect 23954 -780 23966 -720
rect 24000 -780 24012 -720
rect 23954 -792 24012 -780
rect 24084 -720 24142 -708
rect 24084 -780 24096 -720
rect 24130 -780 24142 -720
rect 24084 -792 24142 -780
rect 24172 -720 24230 -708
rect 24172 -780 24184 -720
rect 24218 -780 24230 -720
rect 69466 -720 69524 -708
rect 24172 -792 24230 -780
rect 67024 -746 67082 -734
rect 21730 -818 21788 -806
rect 67024 -806 67036 -746
rect 67070 -806 67082 -746
rect 67024 -818 67082 -806
rect 67112 -746 67170 -734
rect 67112 -806 67124 -746
rect 67158 -806 67170 -746
rect 67112 -818 67170 -806
rect 67242 -746 67300 -734
rect 67242 -806 67254 -746
rect 67288 -806 67300 -746
rect 67242 -818 67300 -806
rect 67330 -746 67388 -734
rect 67330 -806 67342 -746
rect 67376 -806 67388 -746
rect 69466 -780 69478 -720
rect 69512 -780 69524 -720
rect 69466 -792 69524 -780
rect 69554 -720 69612 -708
rect 69554 -780 69566 -720
rect 69600 -780 69612 -720
rect 69554 -792 69612 -780
rect 69684 -720 69742 -708
rect 69684 -780 69696 -720
rect 69730 -780 69742 -720
rect 69684 -792 69742 -780
rect 69772 -720 69830 -708
rect 69772 -780 69784 -720
rect 69818 -780 69830 -720
rect 92266 -720 92324 -708
rect 69772 -792 69830 -780
rect 89824 -746 89882 -734
rect 67330 -818 67388 -806
rect 89824 -806 89836 -746
rect 89870 -806 89882 -746
rect 89824 -818 89882 -806
rect 89912 -746 89970 -734
rect 89912 -806 89924 -746
rect 89958 -806 89970 -746
rect 89912 -818 89970 -806
rect 90042 -746 90100 -734
rect 90042 -806 90054 -746
rect 90088 -806 90100 -746
rect 90042 -818 90100 -806
rect 90130 -746 90188 -734
rect 90130 -806 90142 -746
rect 90176 -806 90188 -746
rect 92266 -780 92278 -720
rect 92312 -780 92324 -720
rect 92266 -792 92324 -780
rect 92354 -720 92412 -708
rect 92354 -780 92366 -720
rect 92400 -780 92412 -720
rect 92354 -792 92412 -780
rect 92484 -720 92542 -708
rect 92484 -780 92496 -720
rect 92530 -780 92542 -720
rect 92484 -792 92542 -780
rect 92572 -720 92630 -708
rect 92572 -780 92584 -720
rect 92618 -780 92630 -720
rect 92572 -792 92630 -780
rect 90130 -818 90188 -806
<< pdiff >>
rect 23866 -338 23924 -326
rect 21424 -364 21482 -352
rect 21424 -592 21436 -364
rect 21470 -592 21482 -364
rect 21424 -604 21482 -592
rect 21512 -364 21570 -352
rect 21512 -592 21524 -364
rect 21558 -592 21570 -364
rect 21512 -604 21570 -592
rect 21642 -364 21700 -352
rect 21642 -592 21654 -364
rect 21688 -592 21700 -364
rect 21642 -604 21700 -592
rect 21730 -364 21788 -352
rect 21730 -592 21742 -364
rect 21776 -592 21788 -364
rect 23866 -566 23878 -338
rect 23912 -566 23924 -338
rect 23866 -578 23924 -566
rect 23954 -338 24012 -326
rect 23954 -566 23966 -338
rect 24000 -566 24012 -338
rect 23954 -578 24012 -566
rect 24084 -338 24142 -326
rect 24084 -566 24096 -338
rect 24130 -566 24142 -338
rect 24084 -578 24142 -566
rect 24172 -338 24230 -326
rect 24172 -566 24184 -338
rect 24218 -566 24230 -338
rect 69466 -338 69524 -326
rect 24172 -578 24230 -566
rect 67024 -364 67082 -352
rect 21730 -604 21788 -592
rect 67024 -592 67036 -364
rect 67070 -592 67082 -364
rect 67024 -604 67082 -592
rect 67112 -364 67170 -352
rect 67112 -592 67124 -364
rect 67158 -592 67170 -364
rect 67112 -604 67170 -592
rect 67242 -364 67300 -352
rect 67242 -592 67254 -364
rect 67288 -592 67300 -364
rect 67242 -604 67300 -592
rect 67330 -364 67388 -352
rect 67330 -592 67342 -364
rect 67376 -592 67388 -364
rect 69466 -566 69478 -338
rect 69512 -566 69524 -338
rect 69466 -578 69524 -566
rect 69554 -338 69612 -326
rect 69554 -566 69566 -338
rect 69600 -566 69612 -338
rect 69554 -578 69612 -566
rect 69684 -338 69742 -326
rect 69684 -566 69696 -338
rect 69730 -566 69742 -338
rect 69684 -578 69742 -566
rect 69772 -338 69830 -326
rect 69772 -566 69784 -338
rect 69818 -566 69830 -338
rect 92266 -338 92324 -326
rect 69772 -578 69830 -566
rect 89824 -364 89882 -352
rect 67330 -604 67388 -592
rect 89824 -592 89836 -364
rect 89870 -592 89882 -364
rect 89824 -604 89882 -592
rect 89912 -364 89970 -352
rect 89912 -592 89924 -364
rect 89958 -592 89970 -364
rect 89912 -604 89970 -592
rect 90042 -364 90100 -352
rect 90042 -592 90054 -364
rect 90088 -592 90100 -364
rect 90042 -604 90100 -592
rect 90130 -364 90188 -352
rect 90130 -592 90142 -364
rect 90176 -592 90188 -364
rect 92266 -566 92278 -338
rect 92312 -566 92324 -338
rect 92266 -578 92324 -566
rect 92354 -338 92412 -326
rect 92354 -566 92366 -338
rect 92400 -566 92412 -338
rect 92354 -578 92412 -566
rect 92484 -338 92542 -326
rect 92484 -566 92496 -338
rect 92530 -566 92542 -338
rect 92484 -578 92542 -566
rect 92572 -338 92630 -326
rect 92572 -566 92584 -338
rect 92618 -566 92630 -338
rect 92572 -578 92630 -566
rect 90130 -604 90188 -592
<< ndiffc >>
rect 21436 -806 21470 -746
rect 21524 -806 21558 -746
rect 21654 -806 21688 -746
rect 21742 -806 21776 -746
rect 23878 -780 23912 -720
rect 23966 -780 24000 -720
rect 24096 -780 24130 -720
rect 24184 -780 24218 -720
rect 67036 -806 67070 -746
rect 67124 -806 67158 -746
rect 67254 -806 67288 -746
rect 67342 -806 67376 -746
rect 69478 -780 69512 -720
rect 69566 -780 69600 -720
rect 69696 -780 69730 -720
rect 69784 -780 69818 -720
rect 89836 -806 89870 -746
rect 89924 -806 89958 -746
rect 90054 -806 90088 -746
rect 90142 -806 90176 -746
rect 92278 -780 92312 -720
rect 92366 -780 92400 -720
rect 92496 -780 92530 -720
rect 92584 -780 92618 -720
<< pdiffc >>
rect 21436 -592 21470 -364
rect 21524 -592 21558 -364
rect 21654 -592 21688 -364
rect 21742 -592 21776 -364
rect 23878 -566 23912 -338
rect 23966 -566 24000 -338
rect 24096 -566 24130 -338
rect 24184 -566 24218 -338
rect 67036 -592 67070 -364
rect 67124 -592 67158 -364
rect 67254 -592 67288 -364
rect 67342 -592 67376 -364
rect 69478 -566 69512 -338
rect 69566 -566 69600 -338
rect 69696 -566 69730 -338
rect 69784 -566 69818 -338
rect 89836 -592 89870 -364
rect 89924 -592 89958 -364
rect 90054 -592 90088 -364
rect 90142 -592 90176 -364
rect 92278 -566 92312 -338
rect 92366 -566 92400 -338
rect 92496 -566 92530 -338
rect 92584 -566 92618 -338
<< poly >>
rect 23924 -326 23954 -300
rect 24142 -326 24172 -300
rect 69524 -326 69554 -300
rect 69742 -326 69772 -300
rect 92324 -326 92354 -300
rect 92542 -326 92572 -300
rect 21482 -352 21512 -326
rect 21700 -352 21730 -326
rect 67082 -352 67112 -326
rect 67300 -352 67330 -326
rect 21164 -660 21396 -644
rect 21164 -700 21182 -660
rect 21376 -662 21396 -660
rect 21482 -662 21512 -604
rect 21700 -642 21730 -604
rect 21376 -694 21512 -662
rect 21376 -700 21396 -694
rect 21164 -716 21396 -700
rect 21482 -734 21512 -694
rect 21554 -652 21730 -642
rect 21554 -688 21578 -652
rect 21680 -688 21730 -652
rect 21554 -698 21730 -688
rect 23606 -634 23838 -618
rect 23606 -674 23624 -634
rect 23818 -636 23838 -634
rect 23924 -636 23954 -578
rect 24142 -616 24172 -578
rect 89882 -352 89912 -326
rect 90100 -352 90130 -326
rect 23818 -668 23954 -636
rect 23818 -674 23838 -668
rect 23606 -690 23838 -674
rect 21700 -734 21730 -698
rect 23924 -708 23954 -668
rect 23996 -626 24172 -616
rect 23996 -662 24020 -626
rect 24122 -662 24172 -626
rect 23996 -672 24172 -662
rect 24142 -708 24172 -672
rect 66764 -660 66996 -644
rect 66764 -700 66782 -660
rect 66976 -662 66996 -660
rect 67082 -662 67112 -604
rect 67300 -642 67330 -604
rect 66976 -694 67112 -662
rect 66976 -700 66996 -694
rect 66764 -716 66996 -700
rect 67082 -734 67112 -694
rect 67154 -652 67330 -642
rect 67154 -688 67178 -652
rect 67280 -688 67330 -652
rect 67154 -698 67330 -688
rect 69206 -634 69438 -618
rect 69206 -674 69224 -634
rect 69418 -636 69438 -634
rect 69524 -636 69554 -578
rect 69742 -616 69772 -578
rect 69418 -668 69554 -636
rect 69418 -674 69438 -668
rect 69206 -690 69438 -674
rect 67300 -734 67330 -698
rect 69524 -708 69554 -668
rect 69596 -626 69772 -616
rect 69596 -662 69620 -626
rect 69722 -662 69772 -626
rect 69596 -672 69772 -662
rect 69742 -708 69772 -672
rect 89564 -660 89796 -644
rect 89564 -700 89582 -660
rect 89776 -662 89796 -660
rect 89882 -662 89912 -604
rect 90100 -642 90130 -604
rect 89776 -694 89912 -662
rect 89776 -700 89796 -694
rect 23924 -818 23954 -792
rect 24142 -818 24172 -792
rect 89564 -716 89796 -700
rect 89882 -734 89912 -694
rect 89954 -652 90130 -642
rect 89954 -688 89978 -652
rect 90080 -688 90130 -652
rect 89954 -698 90130 -688
rect 92006 -634 92238 -618
rect 92006 -674 92024 -634
rect 92218 -636 92238 -634
rect 92324 -636 92354 -578
rect 92542 -616 92572 -578
rect 92218 -668 92354 -636
rect 92218 -674 92238 -668
rect 92006 -690 92238 -674
rect 90100 -734 90130 -698
rect 92324 -708 92354 -668
rect 92396 -626 92572 -616
rect 92396 -662 92420 -626
rect 92522 -662 92572 -626
rect 92396 -672 92572 -662
rect 92542 -708 92572 -672
rect 69524 -818 69554 -792
rect 69742 -818 69772 -792
rect 92324 -818 92354 -792
rect 92542 -818 92572 -792
rect 21482 -844 21512 -818
rect 21700 -844 21730 -818
rect 67082 -844 67112 -818
rect 67300 -844 67330 -818
rect 89882 -844 89912 -818
rect 90100 -844 90130 -818
<< polycont >>
rect 21182 -700 21376 -660
rect 21578 -688 21680 -652
rect 23624 -674 23818 -634
rect 24020 -662 24122 -626
rect 66782 -700 66976 -660
rect 67178 -688 67280 -652
rect 69224 -674 69418 -634
rect 69620 -662 69722 -626
rect 89582 -700 89776 -660
rect 89978 -688 90080 -652
rect 92024 -674 92218 -634
rect 92420 -662 92522 -626
<< locali >>
rect 23878 -338 23912 -322
rect 21436 -364 21470 -348
rect 21436 -608 21470 -592
rect 21524 -364 21558 -348
rect 21524 -608 21558 -592
rect 21654 -364 21688 -348
rect 21654 -608 21688 -592
rect 21742 -364 21776 -348
rect 23878 -582 23912 -566
rect 23966 -338 24000 -322
rect 23966 -582 24000 -566
rect 24096 -338 24130 -322
rect 24096 -582 24130 -566
rect 24184 -338 24218 -322
rect 69478 -338 69512 -322
rect 24184 -582 24218 -566
rect 67036 -364 67070 -348
rect 21742 -608 21776 -592
rect 67036 -608 67070 -592
rect 67124 -364 67158 -348
rect 67124 -608 67158 -592
rect 67254 -364 67288 -348
rect 67254 -608 67288 -592
rect 67342 -364 67376 -348
rect 69478 -582 69512 -566
rect 69566 -338 69600 -322
rect 69566 -582 69600 -566
rect 69696 -338 69730 -322
rect 69696 -582 69730 -566
rect 69784 -338 69818 -322
rect 92278 -338 92312 -322
rect 69784 -582 69818 -566
rect 89836 -364 89870 -348
rect 67342 -608 67376 -592
rect 89836 -608 89870 -592
rect 89924 -364 89958 -348
rect 89924 -608 89958 -592
rect 90054 -364 90088 -348
rect 90054 -608 90088 -592
rect 90142 -364 90176 -348
rect 92278 -582 92312 -566
rect 92366 -338 92400 -322
rect 92366 -582 92400 -566
rect 92496 -338 92530 -322
rect 92496 -582 92530 -566
rect 92584 -338 92618 -322
rect 92584 -582 92618 -566
rect 90142 -608 90176 -592
rect 23606 -634 23838 -618
rect 21164 -660 21396 -644
rect 21164 -700 21182 -660
rect 21376 -700 21396 -660
rect 21554 -652 21712 -642
rect 21554 -688 21578 -652
rect 21680 -688 21712 -652
rect 21554 -696 21712 -688
rect 23606 -674 23624 -634
rect 23818 -674 23838 -634
rect 23996 -626 24154 -616
rect 23996 -662 24020 -626
rect 24122 -662 24154 -626
rect 69206 -634 69438 -618
rect 23996 -670 24154 -662
rect 66764 -660 66996 -644
rect 23606 -690 23838 -674
rect 21164 -716 21396 -700
rect 66764 -700 66782 -660
rect 66976 -700 66996 -660
rect 67154 -652 67312 -642
rect 67154 -688 67178 -652
rect 67280 -688 67312 -652
rect 67154 -696 67312 -688
rect 69206 -674 69224 -634
rect 69418 -674 69438 -634
rect 69596 -626 69754 -616
rect 69596 -662 69620 -626
rect 69722 -662 69754 -626
rect 92006 -634 92238 -618
rect 69596 -670 69754 -662
rect 89564 -660 89796 -644
rect 69206 -690 69438 -674
rect 23878 -720 23912 -704
rect 21436 -746 21470 -730
rect 21436 -822 21470 -806
rect 21524 -746 21558 -730
rect 21524 -822 21558 -806
rect 21654 -746 21688 -730
rect 21654 -822 21688 -806
rect 21742 -746 21776 -730
rect 23878 -796 23912 -780
rect 23966 -720 24000 -704
rect 23966 -796 24000 -780
rect 24096 -720 24130 -704
rect 24096 -796 24130 -780
rect 24184 -720 24218 -704
rect 66764 -716 66996 -700
rect 89564 -700 89582 -660
rect 89776 -700 89796 -660
rect 89954 -652 90112 -642
rect 89954 -688 89978 -652
rect 90080 -688 90112 -652
rect 89954 -696 90112 -688
rect 92006 -674 92024 -634
rect 92218 -674 92238 -634
rect 92396 -626 92554 -616
rect 92396 -662 92420 -626
rect 92522 -662 92554 -626
rect 92396 -670 92554 -662
rect 92006 -690 92238 -674
rect 69478 -720 69512 -704
rect 24184 -796 24218 -780
rect 67036 -746 67070 -730
rect 21742 -822 21776 -806
rect 67036 -822 67070 -806
rect 67124 -746 67158 -730
rect 67124 -822 67158 -806
rect 67254 -746 67288 -730
rect 67254 -822 67288 -806
rect 67342 -746 67376 -730
rect 69478 -796 69512 -780
rect 69566 -720 69600 -704
rect 69566 -796 69600 -780
rect 69696 -720 69730 -704
rect 69696 -796 69730 -780
rect 69784 -720 69818 -704
rect 89564 -716 89796 -700
rect 92278 -720 92312 -704
rect 69784 -796 69818 -780
rect 89836 -746 89870 -730
rect 67342 -822 67376 -806
rect 89836 -822 89870 -806
rect 89924 -746 89958 -730
rect 89924 -822 89958 -806
rect 90054 -746 90088 -730
rect 90054 -822 90088 -806
rect 90142 -746 90176 -730
rect 92278 -796 92312 -780
rect 92366 -720 92400 -704
rect 92366 -796 92400 -780
rect 92496 -720 92530 -704
rect 92496 -796 92530 -780
rect 92584 -720 92618 -704
rect 92584 -796 92618 -780
rect 90142 -822 90176 -806
<< viali >>
rect 21436 -592 21470 -364
rect 21524 -592 21558 -364
rect 21654 -592 21688 -364
rect 21742 -592 21776 -364
rect 23878 -566 23912 -338
rect 23966 -566 24000 -338
rect 24096 -566 24130 -338
rect 24184 -566 24218 -338
rect 67036 -592 67070 -364
rect 67124 -592 67158 -364
rect 67254 -592 67288 -364
rect 67342 -592 67376 -364
rect 69478 -566 69512 -338
rect 69566 -566 69600 -338
rect 69696 -566 69730 -338
rect 69784 -566 69818 -338
rect 89836 -592 89870 -364
rect 89924 -592 89958 -364
rect 90054 -592 90088 -364
rect 90142 -592 90176 -364
rect 92278 -566 92312 -338
rect 92366 -566 92400 -338
rect 92496 -566 92530 -338
rect 92584 -566 92618 -338
rect 21182 -700 21376 -660
rect 21578 -688 21680 -652
rect 23624 -674 23818 -634
rect 24020 -662 24122 -626
rect 66782 -700 66976 -660
rect 67178 -688 67280 -652
rect 69224 -674 69418 -634
rect 69620 -662 69722 -626
rect 21436 -806 21470 -746
rect 21524 -806 21558 -746
rect 21654 -806 21688 -746
rect 21742 -806 21776 -746
rect 23878 -780 23912 -720
rect 23966 -780 24000 -720
rect 24096 -780 24130 -720
rect 89582 -700 89776 -660
rect 89978 -688 90080 -652
rect 92024 -674 92218 -634
rect 92420 -662 92522 -626
rect 24184 -780 24218 -720
rect 67036 -806 67070 -746
rect 67124 -806 67158 -746
rect 67254 -806 67288 -746
rect 67342 -806 67376 -746
rect 69478 -780 69512 -720
rect 69566 -780 69600 -720
rect 69696 -780 69730 -720
rect 69784 -780 69818 -720
rect 89836 -806 89870 -746
rect 89924 -806 89958 -746
rect 90054 -806 90088 -746
rect 90142 -806 90176 -746
rect 92278 -780 92312 -720
rect 92366 -780 92400 -720
rect 92496 -780 92530 -720
rect 92584 -780 92618 -720
<< metal1 >>
rect 42772 2324 45564 2464
rect 42772 2032 42856 2324
rect 45466 2032 45564 2324
rect 42772 1920 45564 2032
rect 19111 246 22847 265
rect 18528 108 22847 246
rect 18528 -688 18660 108
rect 19660 51 22847 108
rect 19660 -688 19866 51
rect 22633 -86 22847 51
rect 44248 18 44824 1920
rect 64751 753 68407 1051
rect 21424 -286 24134 -86
rect 43424 -286 46134 18
rect 64795 -40 65093 753
rect 67024 -2 67352 18
rect 68109 -2 68407 753
rect 85356 422 85882 546
rect 68578 -2 69734 18
rect 64022 -158 65968 -40
rect 21424 -300 23750 -286
rect 21436 -304 21689 -300
rect 21436 -352 21470 -304
rect 21654 -352 21688 -304
rect 23878 -326 23912 -286
rect 24096 -326 24130 -286
rect 43424 -300 45750 -286
rect 23872 -338 23918 -326
rect 21430 -364 21476 -352
rect 21430 -592 21436 -364
rect 21470 -592 21476 -364
rect 21430 -604 21476 -592
rect 21518 -364 21564 -352
rect 21518 -592 21524 -364
rect 21558 -592 21564 -364
rect 21518 -604 21564 -592
rect 21648 -364 21694 -352
rect 21648 -592 21654 -364
rect 21688 -592 21694 -364
rect 21648 -604 21694 -592
rect 21736 -364 21782 -352
rect 21736 -592 21742 -364
rect 21776 -572 21782 -364
rect 23872 -566 23878 -338
rect 23912 -566 23918 -338
rect 21776 -592 21784 -572
rect 23872 -578 23918 -566
rect 23960 -338 24006 -326
rect 23960 -566 23966 -338
rect 24000 -566 24006 -338
rect 23960 -578 24006 -566
rect 24090 -338 24136 -326
rect 24090 -566 24096 -338
rect 24130 -566 24136 -338
rect 24090 -578 24136 -566
rect 24178 -338 24224 -326
rect 24178 -566 24184 -338
rect 24218 -566 24224 -338
rect 24178 -578 24224 -566
rect 64022 -568 64246 -158
rect 65726 -568 65968 -158
rect 67024 -286 69734 -2
rect 67024 -300 69350 -286
rect 67036 -304 67289 -300
rect 67036 -352 67070 -304
rect 67254 -352 67288 -304
rect 69478 -326 69512 -286
rect 69696 -326 69730 -286
rect 69472 -338 69518 -326
rect 21736 -604 21784 -592
rect 21524 -642 21558 -604
rect 21740 -614 21784 -604
rect 21740 -618 23726 -614
rect 23966 -616 24000 -578
rect 21740 -626 23838 -618
rect 21740 -630 23624 -626
rect 18528 -798 19866 -688
rect 21164 -652 21396 -644
rect 21164 -710 21182 -652
rect 21376 -710 21396 -652
rect 21164 -716 21396 -710
rect 21524 -652 21712 -642
rect 21524 -688 21578 -652
rect 21680 -688 21712 -652
rect 21524 -698 21712 -688
rect 21742 -684 23624 -630
rect 23818 -684 23838 -626
rect 21742 -690 23838 -684
rect 23966 -626 24154 -616
rect 23966 -662 24020 -626
rect 24122 -662 24154 -626
rect 23966 -672 24154 -662
rect 24184 -638 24218 -578
rect 43740 -614 43784 -572
rect 43740 -630 45726 -614
rect 43760 -634 45726 -630
rect 24184 -666 24470 -638
rect 21742 -692 23726 -690
rect 21524 -734 21558 -698
rect 21742 -734 21776 -692
rect 23966 -708 24000 -672
rect 24184 -708 24218 -666
rect 23872 -720 23918 -708
rect 21430 -746 21476 -734
rect 19111 -957 19325 -798
rect 21430 -806 21436 -746
rect 21470 -806 21476 -746
rect 21430 -818 21476 -806
rect 21518 -746 21564 -734
rect 21518 -806 21524 -746
rect 21558 -806 21564 -746
rect 21518 -818 21564 -806
rect 21648 -746 21694 -734
rect 21648 -806 21654 -746
rect 21688 -806 21694 -746
rect 21648 -818 21694 -806
rect 21736 -746 21782 -734
rect 21736 -806 21742 -746
rect 21776 -806 21782 -746
rect 23872 -780 23878 -720
rect 23912 -780 23918 -720
rect 23872 -792 23918 -780
rect 23960 -720 24006 -708
rect 23960 -780 23966 -720
rect 24000 -780 24006 -720
rect 23960 -792 24006 -780
rect 24090 -720 24136 -708
rect 24090 -780 24096 -720
rect 24130 -780 24136 -720
rect 24090 -792 24136 -780
rect 24178 -720 24224 -708
rect 24178 -780 24184 -720
rect 24218 -780 24224 -720
rect 24178 -792 24224 -780
rect 21736 -818 21782 -806
rect 21436 -919 21470 -818
rect 21654 -919 21688 -818
rect 22646 -919 22974 -914
rect 23878 -919 23912 -792
rect 24096 -820 24135 -792
rect 24101 -919 24135 -820
rect 21436 -953 24135 -919
rect 22646 -1438 22974 -953
rect 24442 -986 24470 -666
rect 43754 -692 45726 -634
rect 46244 -666 46470 -638
rect 64022 -662 65968 -568
rect 67030 -364 67076 -352
rect 67030 -592 67036 -364
rect 67070 -592 67076 -364
rect 67030 -604 67076 -592
rect 67118 -364 67164 -352
rect 67118 -592 67124 -364
rect 67158 -592 67164 -364
rect 67118 -604 67164 -592
rect 67248 -364 67294 -352
rect 67248 -592 67254 -364
rect 67288 -592 67294 -364
rect 67248 -604 67294 -592
rect 67336 -364 67382 -352
rect 67336 -592 67342 -364
rect 67376 -572 67382 -364
rect 69472 -566 69478 -338
rect 69512 -566 69518 -338
rect 67376 -592 67384 -572
rect 69472 -578 69518 -566
rect 69560 -338 69606 -326
rect 69560 -566 69566 -338
rect 69600 -566 69606 -338
rect 69560 -578 69606 -566
rect 69690 -338 69736 -326
rect 69690 -566 69696 -338
rect 69730 -566 69736 -338
rect 69690 -578 69736 -566
rect 69778 -338 69824 -326
rect 69778 -566 69784 -338
rect 69818 -566 69824 -338
rect 69778 -578 69824 -566
rect 85356 -466 85468 422
rect 85748 18 85882 422
rect 90648 18 91224 84
rect 85748 -286 92534 18
rect 85748 -300 92150 -286
rect 85748 -466 85882 -300
rect 89836 -304 90089 -300
rect 89836 -352 89870 -304
rect 90054 -352 90088 -304
rect 92278 -326 92312 -286
rect 92496 -326 92530 -286
rect 92272 -338 92318 -326
rect 67336 -604 67384 -592
rect 67124 -642 67158 -604
rect 67340 -614 67384 -604
rect 67340 -618 69326 -614
rect 69566 -616 69600 -578
rect 67340 -626 69438 -618
rect 67340 -630 69224 -626
rect 66764 -652 66996 -644
rect 43436 -919 43470 -812
rect 43654 -919 43688 -812
rect 44646 -919 44974 -914
rect 45878 -919 45912 -786
rect 46101 -919 46135 -773
rect 43436 -953 46135 -919
rect 24438 -1008 24916 -986
rect 24438 -1128 24454 -1008
rect 24892 -1128 24916 -1008
rect 24438 -1148 24916 -1128
rect 24442 -1154 24470 -1148
rect 21842 -1530 24278 -1438
rect 44646 -1484 44974 -953
rect 46442 -986 46470 -666
rect 66764 -710 66782 -652
rect 66976 -710 66996 -652
rect 66764 -716 66996 -710
rect 67124 -652 67312 -642
rect 67124 -688 67178 -652
rect 67280 -688 67312 -652
rect 67124 -698 67312 -688
rect 67342 -684 69224 -630
rect 69418 -684 69438 -626
rect 67342 -690 69438 -684
rect 69566 -626 69754 -616
rect 69566 -662 69620 -626
rect 69722 -662 69754 -626
rect 69566 -672 69754 -662
rect 69784 -638 69818 -578
rect 85356 -606 85882 -466
rect 89830 -364 89876 -352
rect 89830 -592 89836 -364
rect 89870 -592 89876 -364
rect 89830 -604 89876 -592
rect 89918 -364 89964 -352
rect 89918 -592 89924 -364
rect 89958 -592 89964 -364
rect 89918 -604 89964 -592
rect 90048 -364 90094 -352
rect 90048 -592 90054 -364
rect 90088 -592 90094 -364
rect 90048 -604 90094 -592
rect 90136 -364 90182 -352
rect 90136 -592 90142 -364
rect 90176 -572 90182 -364
rect 92272 -566 92278 -338
rect 92312 -566 92318 -338
rect 90176 -592 90184 -572
rect 92272 -578 92318 -566
rect 92360 -338 92406 -326
rect 92360 -566 92366 -338
rect 92400 -566 92406 -338
rect 92360 -578 92406 -566
rect 92490 -338 92536 -326
rect 92490 -566 92496 -338
rect 92530 -566 92536 -338
rect 92490 -578 92536 -566
rect 92578 -338 92624 -326
rect 92578 -566 92584 -338
rect 92618 -566 92624 -338
rect 92578 -578 92624 -566
rect 90136 -604 90184 -592
rect 69784 -666 70070 -638
rect 89924 -642 89958 -604
rect 90140 -614 90184 -604
rect 90140 -618 92126 -614
rect 92366 -616 92400 -578
rect 90140 -626 92238 -618
rect 90140 -630 92024 -626
rect 67342 -692 69326 -690
rect 67124 -734 67158 -698
rect 67342 -734 67376 -692
rect 69566 -708 69600 -672
rect 69784 -708 69818 -666
rect 69472 -720 69518 -708
rect 67030 -746 67076 -734
rect 67030 -806 67036 -746
rect 67070 -806 67076 -746
rect 67030 -818 67076 -806
rect 67118 -746 67164 -734
rect 67118 -806 67124 -746
rect 67158 -806 67164 -746
rect 67118 -818 67164 -806
rect 67248 -746 67294 -734
rect 67248 -806 67254 -746
rect 67288 -806 67294 -746
rect 67248 -818 67294 -806
rect 67336 -746 67382 -734
rect 67336 -806 67342 -746
rect 67376 -806 67382 -746
rect 69472 -780 69478 -720
rect 69512 -780 69518 -720
rect 69472 -792 69518 -780
rect 69560 -720 69606 -708
rect 69560 -780 69566 -720
rect 69600 -780 69606 -720
rect 69560 -792 69606 -780
rect 69690 -720 69736 -708
rect 69690 -780 69696 -720
rect 69730 -780 69736 -720
rect 69690 -792 69736 -780
rect 69778 -720 69824 -708
rect 69778 -780 69784 -720
rect 69818 -780 69824 -720
rect 69778 -792 69824 -780
rect 67336 -818 67382 -806
rect 67036 -937 67070 -818
rect 67254 -937 67288 -818
rect 69478 -937 69512 -792
rect 69696 -937 69730 -792
rect 67036 -963 69730 -937
rect 67036 -971 69723 -963
rect 46438 -1008 46916 -986
rect 46438 -1128 46454 -1008
rect 46892 -1128 46916 -1008
rect 46438 -1148 46916 -1128
rect 46442 -1154 46470 -1148
rect 21842 -2010 21962 -1530
rect 24086 -2010 24278 -1530
rect 21842 -2100 24278 -2010
rect 43742 -1598 45968 -1484
rect 43742 -2074 43874 -1598
rect 45832 -2074 45968 -1598
rect 22646 -2102 22974 -2100
rect 43742 -2130 45968 -2074
rect 68006 -1496 68720 -971
rect 70042 -982 70070 -666
rect 89564 -652 89796 -644
rect 89564 -710 89582 -652
rect 89776 -710 89796 -652
rect 89564 -716 89796 -710
rect 89924 -652 90112 -642
rect 89924 -688 89978 -652
rect 90080 -688 90112 -652
rect 89924 -698 90112 -688
rect 90142 -684 92024 -630
rect 92218 -684 92238 -626
rect 90142 -690 92238 -684
rect 92366 -626 92554 -616
rect 92366 -662 92420 -626
rect 92522 -662 92554 -626
rect 92366 -672 92554 -662
rect 92584 -638 92618 -578
rect 92584 -666 92870 -638
rect 90142 -692 92126 -690
rect 89924 -734 89958 -698
rect 90142 -734 90176 -692
rect 92366 -708 92400 -672
rect 92584 -708 92618 -666
rect 92272 -720 92318 -708
rect 89830 -746 89876 -734
rect 89830 -806 89836 -746
rect 89870 -806 89876 -746
rect 89830 -818 89876 -806
rect 89918 -746 89964 -734
rect 89918 -806 89924 -746
rect 89958 -806 89964 -746
rect 89918 -818 89964 -806
rect 90048 -746 90094 -734
rect 90048 -806 90054 -746
rect 90088 -806 90094 -746
rect 90048 -818 90094 -806
rect 90136 -746 90182 -734
rect 90136 -806 90142 -746
rect 90176 -806 90182 -746
rect 92272 -780 92278 -720
rect 92312 -780 92318 -720
rect 92272 -792 92318 -780
rect 92360 -720 92406 -708
rect 92360 -780 92366 -720
rect 92400 -780 92406 -720
rect 92360 -792 92406 -780
rect 92490 -720 92536 -708
rect 92490 -780 92496 -720
rect 92530 -780 92536 -720
rect 92490 -792 92536 -780
rect 92578 -720 92624 -708
rect 92578 -780 92584 -720
rect 92618 -780 92624 -720
rect 92578 -792 92624 -780
rect 90136 -818 90182 -806
rect 70008 -1000 70554 -982
rect 70008 -1142 70054 -1000
rect 70486 -1008 70554 -1000
rect 70492 -1128 70554 -1008
rect 89836 -1003 89870 -818
rect 90054 -1003 90088 -818
rect 90806 -1003 91430 -1002
rect 92278 -1003 92312 -792
rect 92496 -1003 92530 -792
rect 92842 -986 92870 -666
rect 89836 -1037 92530 -1003
rect 92838 -988 93316 -986
rect 92838 -1024 93564 -988
rect 70486 -1142 70554 -1128
rect 70008 -1148 70554 -1142
rect 70042 -1154 70070 -1148
rect 68006 -2038 68072 -1496
rect 68668 -2038 68720 -1496
rect 68006 -2108 68720 -2038
rect 90806 -1516 91430 -1037
rect 92838 -1102 92884 -1024
rect 93526 -1102 93564 -1024
rect 92838 -1142 93564 -1102
rect 92838 -1148 93316 -1142
rect 92842 -1154 92870 -1148
rect 90806 -2032 90888 -1516
rect 91352 -2032 91430 -1516
rect 90806 -2100 91430 -2032
<< via1 >>
rect 42856 2032 45466 2324
rect 18660 -688 19660 108
rect 64246 -568 65726 -158
rect 21182 -660 21376 -652
rect 21182 -700 21376 -660
rect 21182 -710 21376 -700
rect 23624 -634 23818 -626
rect 23624 -674 23818 -634
rect 23624 -684 23818 -674
rect 85468 -466 85748 422
rect 24454 -1128 24892 -1008
rect 66782 -660 66976 -652
rect 66782 -700 66976 -660
rect 66782 -710 66976 -700
rect 69224 -634 69418 -626
rect 69224 -674 69418 -634
rect 69224 -684 69418 -674
rect 46454 -1128 46892 -1008
rect 21962 -2010 24086 -1530
rect 43874 -2074 45832 -1598
rect 89582 -660 89776 -652
rect 89582 -700 89776 -660
rect 89582 -710 89776 -700
rect 92024 -634 92218 -626
rect 92024 -674 92218 -634
rect 92024 -684 92218 -674
rect 70054 -1008 70486 -1000
rect 70054 -1128 70492 -1008
rect 70054 -1142 70486 -1128
rect 68072 -2038 68668 -1496
rect 92884 -1102 93526 -1024
rect 90888 -2032 91352 -1516
<< metal2 >>
rect 21150 23582 24582 23700
rect 44708 23612 47926 23696
rect 68102 23628 71614 23698
rect 91594 23618 95064 23686
rect 21188 21502 24620 21620
rect 44694 21526 47912 21610
rect 68088 21572 71600 21606
rect 68088 21536 71674 21572
rect 91596 21540 95066 21608
rect 71468 21496 71674 21536
rect 21158 19414 24590 19532
rect 44680 19444 47898 19528
rect 68092 19460 71604 19530
rect 91586 19452 95056 19520
rect 21102 17328 24640 17440
rect 44708 17362 47926 17446
rect 68002 17382 71514 17452
rect 91608 17366 95078 17434
rect 21090 15320 24628 15374
rect 21090 15254 24634 15320
rect 44688 15278 47906 15362
rect 67996 15292 71508 15362
rect 91594 15282 95064 15350
rect 21096 15224 24634 15254
rect 21100 13288 24638 13320
rect 21062 13238 24638 13288
rect 21090 13224 24638 13238
rect 21090 13156 24628 13224
rect 44740 13192 47958 13276
rect 68014 13206 71526 13276
rect 91650 13196 95120 13264
rect 47894 11194 47974 11258
rect 44722 11172 47974 11194
rect 21068 11062 24606 11158
rect 44722 11110 47940 11172
rect 68010 11116 71522 11186
rect 91648 11108 95118 11176
rect 21024 9100 24594 9106
rect 21024 9030 24610 9100
rect 21024 8962 24594 9030
rect 44742 9020 47960 9104
rect 67982 9034 71494 9104
rect 91658 9030 95128 9098
rect 42772 2324 45564 2464
rect 42772 2032 42856 2324
rect 45466 2032 45564 2324
rect 42772 1920 45564 2032
rect 85356 422 85882 546
rect 18528 108 19866 246
rect 18528 -688 18660 108
rect 19660 -688 19866 108
rect 64022 -158 65968 -40
rect 64022 -568 64246 -158
rect 65726 -568 65968 -158
rect 23606 -626 23838 -618
rect 18528 -798 19866 -688
rect 20856 -652 21396 -644
rect 20856 -710 21182 -652
rect 21376 -710 21396 -652
rect 23606 -684 23624 -626
rect 23818 -684 23838 -626
rect 23606 -690 23838 -684
rect 20856 -716 21396 -710
rect 20856 -726 21226 -716
rect 20856 -1108 20914 -726
rect 21162 -1108 21226 -726
rect 42856 -726 43226 -644
rect 64022 -662 65968 -568
rect 85356 -466 85468 422
rect 85748 -466 85882 422
rect 85356 -606 85882 -466
rect 69206 -626 69438 -618
rect 66456 -652 66996 -644
rect 20856 -1148 21226 -1108
rect 24438 -1008 24916 -986
rect 24438 -1128 24454 -1008
rect 24892 -1128 24916 -1008
rect 24438 -1148 24916 -1128
rect 42856 -1108 42914 -726
rect 43162 -1108 43226 -726
rect 66456 -710 66782 -652
rect 66976 -710 66996 -652
rect 69206 -684 69224 -626
rect 69418 -684 69438 -626
rect 92006 -626 92238 -618
rect 69206 -690 69438 -684
rect 89256 -652 89796 -644
rect 66456 -716 66996 -710
rect 89256 -710 89582 -652
rect 89776 -692 89796 -652
rect 92006 -684 92024 -626
rect 92218 -684 92238 -626
rect 92006 -690 92238 -684
rect 89776 -710 89784 -692
rect 89256 -716 89784 -710
rect 66456 -726 66826 -716
rect 89256 -726 89626 -716
rect 42856 -1148 43226 -1108
rect 46438 -1008 46916 -986
rect 46438 -1128 46454 -1008
rect 46892 -1128 46916 -1008
rect 46438 -1148 46916 -1128
rect 66456 -1108 66514 -726
rect 66762 -1108 66794 -726
rect 66456 -1148 66794 -1108
rect 70038 -1000 70516 -986
rect 70038 -1142 70054 -1000
rect 70486 -1008 70516 -1000
rect 70492 -1128 70516 -1008
rect 70486 -1142 70516 -1128
rect 70038 -1148 70516 -1142
rect 89256 -1108 89314 -726
rect 89562 -1108 89626 -726
rect 89256 -1148 89626 -1108
rect 92844 -1024 93564 -988
rect 92844 -1102 92884 -1024
rect 93526 -1102 93564 -1024
rect 92844 -1142 93564 -1102
rect 21842 -1530 24278 -1438
rect 44457 -1480 44591 -1432
rect 21842 -2010 21962 -1530
rect 24086 -2010 24278 -1530
rect 21842 -2100 24278 -2010
rect 43738 -1598 45966 -1480
rect 43738 -2074 43874 -1598
rect 45834 -2070 45966 -1598
rect 45832 -2074 45966 -2070
rect 43738 -2136 45966 -2074
rect 68006 -1496 68714 -1442
rect 68006 -2038 68072 -1496
rect 68668 -2038 68714 -1496
rect 68006 -2108 68714 -2038
rect 90806 -1516 91436 -1444
rect 90806 -2032 90888 -1516
rect 91352 -2032 91436 -1516
rect 90806 -2100 91436 -2032
<< via2 >>
rect 42856 2032 45466 2324
rect 18660 -688 19660 108
rect 64246 -568 65726 -158
rect 20914 -1108 21162 -726
rect 85468 -466 85748 422
rect 24454 -1128 24892 -1008
rect 42914 -1108 43162 -726
rect 46454 -1128 46892 -1008
rect 66514 -1108 66762 -726
rect 70054 -1142 70486 -1000
rect 89314 -1108 89562 -726
rect 92884 -1102 93526 -1024
rect 21962 -2010 24086 -1530
rect 43882 -2070 45832 -1598
rect 45832 -2070 45834 -1598
rect 68072 -2038 68668 -1496
rect 90888 -2032 91352 -1516
<< metal3 >>
rect 66614 5480 67352 5900
rect 42772 2344 45564 2464
rect 42772 2324 42870 2344
rect 45446 2324 45564 2344
rect 42772 2032 42856 2324
rect 45466 2032 45564 2324
rect 42772 2022 42870 2032
rect 45446 2022 45564 2032
rect 42772 1920 45564 2022
rect 85356 422 85882 546
rect 11256 -984 11420 246
rect 18528 108 19866 246
rect 18528 -688 18660 108
rect 19660 -688 19866 108
rect 18528 -798 19866 -688
rect 20856 -726 21226 -644
rect 20856 -984 20914 -726
rect 11256 -1108 20914 -984
rect 21162 -1108 21226 -726
rect 34772 -908 34984 -600
rect 34776 -984 34984 -908
rect 42856 -726 43226 -644
rect 42856 -984 42914 -726
rect 11256 -1148 21226 -1108
rect 24414 -1008 42914 -984
rect 24414 -1128 24454 -1008
rect 24892 -1108 42914 -1008
rect 43162 -1108 43226 -726
rect 57322 -984 57578 -980
rect 58114 -984 58278 266
rect 64022 -158 65968 -40
rect 64022 -568 64246 -158
rect 65726 -568 65968 -158
rect 64022 -662 65968 -568
rect 85356 -466 85468 422
rect 85748 -466 85882 422
rect 66456 -726 66826 -644
rect 66456 -984 66514 -726
rect 46444 -986 66514 -984
rect 24892 -1128 43226 -1108
rect 24414 -1148 43226 -1128
rect 46438 -1008 66514 -986
rect 46438 -1128 46454 -1008
rect 46892 -1108 66514 -1008
rect 66762 -1108 66826 -726
rect 79584 -984 79766 -974
rect 81768 -984 81840 -596
rect 85356 -606 85882 -466
rect 89256 -726 89626 -644
rect 89256 -984 89314 -726
rect 46892 -1128 66826 -1108
rect 46438 -1148 66826 -1128
rect 69948 -1000 89314 -984
rect 69948 -1142 70054 -1000
rect 70486 -1108 89314 -1000
rect 89562 -984 89626 -726
rect 105264 -984 105428 262
rect 89562 -1108 89636 -984
rect 92844 -986 102348 -984
rect 70486 -1142 89636 -1108
rect 69948 -1148 89636 -1142
rect 92838 -988 102348 -986
rect 102996 -988 105428 -984
rect 92838 -1024 105428 -988
rect 92838 -1102 92884 -1024
rect 93526 -1102 105428 -1024
rect 92838 -1148 105428 -1102
rect 57322 -1154 57578 -1148
rect 21842 -1530 24278 -1438
rect 21842 -1540 21962 -1530
rect 21842 -1992 21958 -1540
rect 21842 -2010 21962 -1992
rect 24086 -2010 24278 -1530
rect 21842 -2100 24278 -2010
rect 43738 -1598 45966 -1480
rect 43738 -2070 43882 -1598
rect 45834 -2070 45966 -1598
rect 43738 -2136 45966 -2070
rect 68006 -1482 68714 -1442
rect 68006 -1496 68086 -1482
rect 68006 -2038 68072 -1496
rect 68006 -2060 68086 -2038
rect 68690 -2060 68714 -1482
rect 68006 -2108 68714 -2060
rect 90806 -1500 91436 -1444
rect 90806 -2022 90874 -1500
rect 91368 -2022 91436 -1500
rect 90806 -2032 90888 -2022
rect 91352 -2032 91436 -2022
rect 90806 -2100 91436 -2032
<< via3 >>
rect 42870 2324 45446 2344
rect 42870 2032 45446 2324
rect 42870 2022 45446 2032
rect 18660 -688 19660 108
rect 64246 -568 65726 -158
rect 85468 -466 85748 422
rect 21958 -1992 21962 -1540
rect 21962 -1992 24056 -1540
rect 43900 -2060 45818 -1610
rect 68086 -1496 68690 -1482
rect 68086 -2038 68668 -1496
rect 68668 -2038 68690 -1496
rect 68086 -2060 68690 -2038
rect 90874 -1516 91368 -1500
rect 90874 -2022 90888 -1516
rect 90888 -2022 91352 -1516
rect 91352 -2022 91368 -1516
<< metal4 >>
rect 148 -405 806 3223
rect 18528 108 19866 246
rect 18528 -405 18660 108
rect 148 -688 18660 -405
rect 19660 -405 19866 108
rect 19660 -688 19873 -405
rect 148 -1063 19873 -688
rect 148 -2965 806 -1063
rect 21820 -1540 24270 -1442
rect 21820 -1992 21958 -1540
rect 24056 -1992 24270 -1540
rect 21820 -2144 24270 -1992
rect 39674 -2965 40246 2490
rect 54140 -26 54791 3155
rect 85338 422 85910 2496
rect 54140 -100 58996 -26
rect 60726 -100 66423 -26
rect 54140 -158 66423 -100
rect 54140 -568 64246 -158
rect 65726 -568 66423 -158
rect 54140 -677 66423 -568
rect 85338 -466 85468 422
rect 85748 -466 85910 422
rect 43740 -1610 45990 -1450
rect 43740 -2060 43900 -1610
rect 45818 -2060 45990 -1610
rect 43740 -2136 45990 -2060
rect 54140 -2965 54791 -677
rect 67934 -1482 68746 -1428
rect 67934 -2060 68086 -1482
rect 68690 -2060 68746 -1482
rect 67934 -2156 68746 -2060
rect 85338 -2965 85910 -466
rect 90812 -1500 91442 -1458
rect 90812 -2022 90874 -1500
rect 91368 -2022 91442 -1500
rect 90812 -2104 91442 -2022
rect 102295 -2965 102953 3073
rect 148 -3623 102953 -2965
rect 39674 -3698 40246 -3623
rect 85338 -3814 85910 -3623
<< via4 >>
rect 21958 -1992 24056 -1540
rect 43900 -2060 45818 -1610
rect 68086 -2060 68690 -1482
rect 90894 -2022 91360 -1506
<< metal5 >>
rect -446 -1444 212 9305
rect 20023 3555 22324 4145
rect 115938 3235 116596 18609
rect 14972 -1444 15708 2994
rect 29098 -1444 29834 2468
rect 32490 1924 33300 3181
rect 61808 -1444 62544 3230
rect 73942 -1444 74678 2760
rect 106759 2577 116596 3235
rect 115938 -1444 116596 2577
rect -446 -1482 116596 -1444
rect -446 -1540 68086 -1482
rect -446 -1963 21958 -1540
rect -444 -1992 21958 -1963
rect 24056 -1610 68086 -1540
rect 24056 -1992 43900 -1610
rect -444 -2060 43900 -1992
rect 45818 -2060 68086 -1610
rect 68690 -1506 116596 -1482
rect 68690 -2022 90894 -1506
rect 91360 -2022 116596 -1506
rect 68690 -2060 116596 -2022
rect -444 -2149 116596 -2060
rect -444 -2180 116410 -2149
use buffer_digital  buffer_digital_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698389822
transform 1 0 43438 0 1 -846
box -274 0 412 576
use buffer_digital  buffer_digital_1
timestamp 1698389822
transform 1 0 45880 0 1 -820
box -274 0 412 576
use charge_pump3  charge_pump3_0
timestamp 1698660782
transform 1 0 22380 0 -1 24868
box 498 -3206 23756 25756
use charge_pump3  charge_pump3_1
timestamp 1698660782
transform 1 0 69294 0 -1 24874
box 498 -3206 23756 25756
use charge_pump  charge_pump_0 ~/Desktop/charge_pumps2/layout_files2
timestamp 1698659501
transform 1 0 -1210 0 1 7820
box 498 -7862 23756 19014
use charge_pump  charge_pump_1
timestamp 1698659501
transform 1 0 45712 0 1 7856
box 498 -7862 23756 19014
use charge_pump  charge_pump_2
timestamp 1698659501
transform 1 0 92840 0 1 7848
box 498 -7862 23756 19014
<< end >>
