magic
tech sky130A
magscale 1 2
timestamp 1727642364
<< nwell >>
rect 7832 -796 8184 -624
rect 7902 -802 8140 -796
<< pwell >>
rect 7804 -1458 8236 -1262
rect 7800 -1626 8240 -1458
<< psubdiff >>
rect 5661 -409 5748 -383
rect 5661 -450 5688 -409
rect 5722 -450 5748 -409
rect 5661 -475 5748 -450
rect 7852 -1498 8188 -1474
rect 7852 -1556 7886 -1498
rect 8162 -1556 8188 -1498
rect 7852 -1584 8188 -1556
<< nsubdiff >>
rect 7912 -686 8128 -660
rect 7912 -722 7946 -686
rect 8094 -722 8128 -686
rect 7912 -750 8128 -722
<< psubdiffcont >>
rect 5688 -450 5722 -409
rect 7886 -1556 8162 -1498
<< nsubdiffcont >>
rect 7946 -722 8094 -686
<< poly >>
rect 38 -356 173 -322
rect 38 -375 72 -356
rect 932 -359 1061 -329
rect 932 -402 962 -359
rect 1890 -362 2013 -332
rect 2848 -352 2977 -322
rect 3830 -329 3860 -324
rect 1890 -394 1920 -362
rect 2848 -384 2878 -352
rect 3830 -359 3959 -329
rect 4772 -356 4901 -326
rect 3830 -386 3860 -359
rect 4772 -388 4802 -356
<< locali >>
rect 302 -290 988 -258
rect 5661 -409 5748 -383
rect 5661 -451 5687 -409
rect 5722 -451 5748 -409
rect 5661 -475 5748 -451
rect -16 -612 5796 -526
rect -16 -614 666 -612
rect 7912 -686 8128 -660
rect 7912 -722 7946 -686
rect 8094 -722 8128 -686
rect 7912 -750 8128 -722
rect 8050 -844 8088 -750
rect 7936 -1474 7986 -1360
rect 7852 -1498 8188 -1474
rect 7852 -1556 7886 -1498
rect 8162 -1556 8188 -1498
rect 7852 -1584 8188 -1556
<< viali >>
rect 5687 -450 5688 -409
rect 5688 -450 5722 -409
rect 5687 -451 5722 -450
<< metal1 >>
rect -224 1564 6008 1598
rect -224 1534 6036 1564
rect -242 1343 -232 1534
rect -274 1330 -232 1343
rect 5994 1425 6036 1534
rect 5994 1383 6295 1425
rect 5994 1330 6036 1383
rect -274 1309 6036 1330
rect -224 1244 6036 1309
rect 424 1064 528 1244
rect 5503 1228 5623 1244
rect 5740 1217 5856 1244
rect 5884 1228 6036 1244
rect -274 960 914 1064
rect -660 465 -344 466
rect -1456 458 -344 465
rect -1456 399 -636 458
rect -2450 -655 -2416 -524
rect -855 -1171 -789 399
rect -660 398 -636 399
rect -374 398 -344 458
rect -660 384 -344 398
rect -274 -578 -170 960
rect 424 930 528 960
rect 2438 884 2524 896
rect 2436 828 2446 884
rect 2508 828 2524 884
rect 2438 824 2524 828
rect 870 244 974 258
rect 870 190 882 244
rect 954 190 974 244
rect 1254 192 1264 250
rect 1346 192 1356 250
rect 2424 192 2434 252
rect 2508 192 2518 252
rect 2812 190 2822 248
rect 2892 190 2902 248
rect 870 188 974 190
rect 5918 -76 6116 -56
rect 5918 -132 5936 -76
rect 6094 -132 6116 -76
rect 5918 -150 6116 -132
rect 6075 -162 6113 -150
rect -12 -432 16 -212
rect 302 -290 988 -264
rect 124 -360 740 -326
rect 882 -420 916 -290
rect 1014 -376 1646 -326
rect 1840 -416 1874 -260
rect 1968 -372 2600 -322
rect -14 -460 790 -432
rect -12 -470 16 -460
rect 878 -472 1680 -420
rect 1840 -454 2646 -416
rect 1844 -468 2646 -454
rect 2794 -424 2828 -260
rect 2934 -372 3560 -330
rect 3780 -424 3814 -266
rect 3920 -376 4546 -334
rect 4722 -420 4756 -274
rect 4854 -374 5480 -332
rect 5680 -397 5728 -213
rect 5680 -409 5730 -397
rect 2794 -476 3596 -424
rect 3778 -476 4580 -424
rect 4720 -472 5522 -420
rect 5680 -451 5687 -409
rect 5722 -451 5730 -409
rect 5680 -464 5730 -451
rect 26 -520 664 -516
rect -16 -526 666 -520
rect -16 -578 5796 -526
rect -274 -612 5796 -578
rect -274 -614 666 -612
rect -274 -682 2 -614
rect -506 -1162 -416 -1160
rect -506 -1171 -190 -1162
rect -855 -1176 -190 -1171
rect -855 -1232 -440 -1176
rect -224 -1232 -190 -1176
rect -855 -1237 -190 -1232
rect -506 -1244 -190 -1237
rect -478 -1246 -190 -1244
rect -924 -1400 -310 -1384
rect -924 -1462 -766 -1400
rect -382 -1462 -310 -1400
rect 826 -1442 836 -1378
rect 926 -1442 936 -1378
rect 1212 -1440 1222 -1376
rect 1312 -1440 1322 -1376
rect 2366 -1386 2480 -1372
rect 2366 -1442 2404 -1386
rect 2472 -1442 2482 -1386
rect 2366 -1444 2480 -1442
rect 2778 -1444 2788 -1390
rect 2852 -1444 2862 -1390
rect -924 -1484 -310 -1462
rect -732 -1516 -700 -1513
rect -804 -1558 -660 -1516
rect -804 -1574 -594 -1558
rect -776 -1588 -594 -1574
rect -776 -1746 -730 -1588
rect -646 -1746 -594 -1588
rect -2480 -1776 -2408 -1764
rect -776 -1796 -594 -1746
rect -170 -1820 5588 -1818
rect 5864 -1820 5962 -178
rect 6253 -825 6295 1383
rect 8232 -1080 8345 -1030
rect 6075 -1120 6113 -1114
rect 6009 -1158 6151 -1120
rect 6009 -1614 6047 -1158
rect 6076 -1204 6166 -1196
rect 6076 -1258 6088 -1204
rect 6148 -1258 6166 -1204
rect 6076 -1276 6166 -1258
rect 6009 -1640 6116 -1614
rect 6009 -1733 6036 -1640
rect 6022 -1758 6036 -1733
rect 6102 -1758 6116 -1640
rect 6022 -1784 6116 -1758
rect -170 -1890 6052 -1820
rect -146 -1936 6052 -1890
rect -154 -1970 -144 -1936
rect -170 -1996 -144 -1970
rect -186 -2114 -144 -1996
rect 6022 -2048 6052 -1936
rect 6278 -2048 6314 -1346
rect 6022 -2084 6314 -2048
rect 6022 -2114 6052 -2084
rect -186 -2162 6052 -2114
rect -146 -2214 6052 -2162
<< via1 >>
rect -232 1330 5994 1534
rect -636 398 -374 458
rect 2446 828 2508 884
rect 882 190 954 244
rect 1264 192 1346 250
rect 2434 192 2508 252
rect 2822 190 2892 248
rect 5936 -132 6094 -76
rect -440 -1232 -224 -1176
rect -766 -1462 -382 -1400
rect 836 -1442 926 -1378
rect 1222 -1440 1312 -1376
rect 2404 -1442 2472 -1386
rect 2788 -1444 2852 -1390
rect -730 -1746 -646 -1588
rect 6088 -1258 6148 -1204
rect 6036 -1758 6102 -1640
rect -144 -2114 6022 -1936
<< metal2 >>
rect -232 1534 5994 1544
rect -232 1320 5994 1330
rect 2438 884 2524 896
rect 2438 828 2446 884
rect 2508 828 2524 884
rect 2438 824 2524 828
rect 2446 818 2508 824
rect -660 458 -344 466
rect -660 398 -636 458
rect -374 398 -344 458
rect -660 384 -344 398
rect -1398 296 1314 326
rect -701 -1286 -671 296
rect 1284 262 1314 296
rect -642 238 -302 246
rect -642 160 -608 238
rect -328 224 -302 238
rect 870 244 974 258
rect 870 224 882 244
rect -328 190 882 224
rect 954 190 974 244
rect 1258 250 1358 262
rect 1258 192 1264 250
rect 1346 192 1358 250
rect 1258 190 1358 192
rect 2434 252 2508 262
rect -328 188 974 190
rect -328 160 -302 188
rect 882 180 954 188
rect 1264 182 1346 190
rect 2434 182 2508 192
rect 2822 248 2892 258
rect 2822 180 2892 190
rect -642 140 -302 160
rect 4746 -80 4874 -70
rect 5918 -76 6116 -56
rect 5918 -132 5936 -76
rect 6094 -132 6116 -76
rect 5918 -150 6116 -132
rect 4746 -166 4874 -156
rect 2764 -732 2872 -722
rect 2764 -808 2872 -798
rect -478 -1176 -190 -1162
rect -478 -1232 -440 -1176
rect -224 -1232 -190 -1176
rect -478 -1246 -190 -1232
rect 6074 -1196 6108 -150
rect 6074 -1204 6166 -1196
rect 6074 -1238 6088 -1204
rect 6076 -1258 6088 -1238
rect 6148 -1258 6166 -1204
rect 6076 -1276 6166 -1258
rect -701 -1316 1284 -1286
rect -700 -1318 1284 -1316
rect -700 -1320 -418 -1318
rect 776 -1366 954 -1364
rect 1252 -1366 1284 -1318
rect 776 -1378 956 -1366
rect -924 -1396 -310 -1384
rect -924 -1460 -768 -1396
rect -382 -1424 -310 -1396
rect 776 -1424 836 -1378
rect -382 -1442 836 -1424
rect 926 -1442 956 -1378
rect -382 -1446 956 -1442
rect 1174 -1376 1334 -1366
rect 1174 -1440 1222 -1376
rect 1312 -1440 1334 -1376
rect 1174 -1446 1334 -1440
rect 2366 -1382 2480 -1372
rect 2366 -1442 2404 -1382
rect 2472 -1442 2480 -1382
rect 2366 -1444 2480 -1442
rect 2788 -1384 2852 -1374
rect -382 -1452 954 -1446
rect 1222 -1450 1312 -1446
rect 2404 -1452 2472 -1444
rect -924 -1462 -766 -1460
rect -382 -1462 -310 -1452
rect 2788 -1454 2852 -1444
rect -924 -1484 -310 -1462
rect -776 -1588 -594 -1558
rect -776 -1746 -730 -1588
rect -646 -1746 -594 -1588
rect 6022 -1640 6116 -1614
rect -776 -1796 -594 -1746
rect 4718 -1712 4846 -1702
rect 6022 -1758 6036 -1640
rect 6102 -1758 6116 -1640
rect 6022 -1784 6116 -1758
rect 4718 -1800 4846 -1790
rect -144 -1936 6022 -1926
rect -144 -2124 6022 -2114
<< via2 >>
rect -232 1330 5994 1534
rect 2446 828 2508 884
rect -636 398 -374 458
rect -608 160 -328 238
rect 2434 192 2508 252
rect 2822 190 2892 248
rect 4746 -156 4874 -80
rect 5936 -132 6094 -76
rect 2764 -798 2872 -732
rect -440 -1232 -224 -1176
rect -768 -1400 -382 -1396
rect -768 -1460 -766 -1400
rect -766 -1460 -382 -1400
rect 2404 -1386 2472 -1382
rect 2404 -1438 2472 -1386
rect 2788 -1390 2852 -1384
rect 2788 -1444 2852 -1390
rect -730 -1746 -646 -1588
rect 4718 -1790 4846 -1712
rect 6036 -1758 6102 -1640
rect -144 -2114 6022 -1936
<< metal3 >>
rect -242 1294 -232 1576
rect 6000 1294 6010 1576
rect 2438 894 2524 896
rect 2430 884 2524 894
rect 2430 866 2446 884
rect 2428 828 2446 866
rect 2508 828 2524 884
rect 2428 824 2524 828
rect 2428 778 2518 824
rect -476 738 -466 744
rect -500 658 -466 738
rect -476 644 -466 658
rect -366 738 -356 744
rect 2428 738 2508 778
rect -366 658 2508 738
rect -366 644 -356 658
rect -660 460 -344 466
rect -660 458 2506 460
rect -660 398 -636 458
rect -374 398 2506 458
rect -660 388 2506 398
rect -660 384 -344 388
rect 2434 274 2506 388
rect 2410 252 2528 274
rect -642 238 -302 246
rect -642 221 -608 238
rect -1130 160 -608 221
rect -328 160 -302 238
rect 2410 192 2434 252
rect 2508 192 2528 252
rect 2410 184 2528 192
rect 2796 248 2914 274
rect 2796 190 2822 248
rect 2892 190 2914 248
rect 2796 184 2914 190
rect -1130 155 -302 160
rect -1130 -1692 -1064 155
rect -642 140 -302 155
rect 2812 -80 2892 184
rect -631 -128 2892 -80
rect 4736 -80 4884 -75
rect -631 -158 2890 -128
rect 4736 -156 4746 -80
rect 4874 -82 4884 -80
rect 5918 -76 6116 -56
rect 5918 -82 5936 -76
rect 4874 -132 5936 -82
rect 6094 -132 6116 -76
rect 4874 -150 6116 -132
rect 4874 -152 6026 -150
rect 4874 -156 4944 -152
rect -631 -1382 -553 -158
rect 4736 -161 4884 -156
rect 2754 -732 2882 -727
rect 2754 -798 2764 -732
rect 2872 -798 2882 -732
rect 2754 -803 2882 -798
rect -470 -988 -460 -890
rect -354 -908 -344 -890
rect 2790 -908 2850 -803
rect -354 -968 2850 -908
rect -354 -988 -344 -968
rect -478 -1173 -190 -1162
rect -478 -1176 2462 -1173
rect -478 -1232 -440 -1176
rect -224 -1232 2462 -1176
rect -478 -1235 2462 -1232
rect -478 -1246 -190 -1235
rect 2400 -1356 2462 -1235
rect 2366 -1382 2482 -1356
rect 2798 -1358 2858 -1356
rect -920 -1396 -308 -1382
rect -920 -1460 -768 -1396
rect -382 -1460 -308 -1396
rect 2366 -1438 2404 -1382
rect 2472 -1438 2482 -1382
rect 2366 -1444 2482 -1438
rect 2772 -1384 2886 -1358
rect 2772 -1444 2788 -1384
rect 2852 -1444 2886 -1384
rect 2772 -1450 2886 -1444
rect -920 -1484 -308 -1460
rect -631 -1485 -553 -1484
rect -1128 -1732 -1064 -1692
rect -776 -1588 -594 -1558
rect -776 -1730 -730 -1588
rect -840 -1732 -730 -1730
rect -1128 -1746 -730 -1732
rect -646 -1730 -594 -1588
rect -646 -1732 -502 -1730
rect 2798 -1732 2858 -1450
rect 6022 -1640 6116 -1614
rect -646 -1746 2858 -1732
rect -1128 -1792 2858 -1746
rect 4708 -1712 4856 -1707
rect 6022 -1712 6036 -1640
rect 4708 -1790 4718 -1712
rect 4846 -1758 6036 -1712
rect 6102 -1758 6116 -1640
rect 4846 -1780 6116 -1758
rect 4846 -1790 4856 -1780
rect 6022 -1784 6116 -1780
rect -1128 -1795 -1064 -1792
rect -776 -1796 -594 -1792
rect 4708 -1795 4856 -1790
rect -154 -1931 6028 -1896
rect -154 -1936 6032 -1931
rect -154 -2114 -144 -1936
rect 6022 -2114 6032 -1936
rect -154 -2119 6032 -2114
<< via3 >>
rect -232 1534 6000 1576
rect -232 1330 5994 1534
rect 5994 1330 6000 1534
rect -232 1294 6000 1330
rect -466 644 -366 744
rect -460 -988 -354 -890
<< metal4 >>
rect -232 1577 6022 1614
rect -233 1576 6022 1577
rect -233 1556 -232 1576
rect -274 1318 -232 1556
rect -233 1294 -232 1318
rect 6000 1294 6022 1576
rect -233 1293 6022 1294
rect -232 1228 6022 1293
rect -232 1214 4944 1228
rect 5714 1214 6022 1228
rect -467 744 -365 745
rect -467 644 -466 744
rect -366 644 -365 744
rect -467 643 -365 644
rect -466 -790 -366 643
rect -466 -890 -352 -790
rect -466 -984 -460 -890
rect -461 -988 -460 -984
rect -354 -984 -352 -890
rect -354 -988 -353 -984
rect -461 -989 -353 -988
use comparator_full_compact  comparator_full_compact_0
timestamp 1698871213
transform 1 0 622 0 1 -292
box -794 -4 5299 1494
use comparator_full_compact  comparator_full_compact_1
timestamp 1698871213
transform 1 0 592 0 1 -1922
box -794 -4 5299 1494
use reference  reference_0
timestamp 1727087973
transform 1 0 -2500 0 1 -1085
box -32 -858 1828 500
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_0
timestamp 1698873245
transform 1 0 389 0 1 -442
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_1
timestamp 1698873245
transform 1 0 1283 0 1 -446
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_2
timestamp 1698873245
transform 1 0 2241 0 1 -444
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_3
timestamp 1698873245
transform 1 0 3199 0 1 -444
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_4
timestamp 1698873245
transform 1 0 4181 0 1 -446
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_5
timestamp 1698873245
transform 1 0 5123 0 1 -446
box -413 -130 413 130
use xnor  xnor_0
timestamp 1727642364
transform 1 0 6222 0 1 -1374
box -147 -48 2062 592
<< labels >>
rlabel metal2 -253 -1302 -253 -1302 1 V+
rlabel via2 -289 -1211 -289 -1211 1 V-
rlabel metal3 -373 430 -373 430 1 V-
rlabel metal2 -369 312 -369 312 1 V+
rlabel via2 -380 200 -380 200 1 Vc+
rlabel metal3 -358 -112 -358 -112 1 Vc-
rlabel metal1 -1384 428 -1384 428 1 V-
rlabel metal2 -692 -1088 -692 -1088 1 V+
port 5 n
rlabel metal4 -418 -746 -418 -746 1 clk
port 9 n
rlabel metal1 -1440 436 -1440 436 1 V-
port 10 n
rlabel metal1 -2430 -558 -2430 -558 1 vdd_ref
rlabel space -2450 -1808 -2450 -1808 1 gnd_ref
<< end >>
