magic
tech sky130A
magscale 1 2
timestamp 1697921677
<< locali >>
rect 2418 3684 4121 3693
rect 2418 3625 4121 3647
rect 2634 3392 2871 3433
rect 3701 3385 3929 3440
rect 2609 2849 2915 2893
rect 3766 2856 4072 2900
rect 2420 2672 4123 2692
rect 4122 2635 4123 2672
rect 2420 2624 4123 2635
<< viali >>
rect 2415 3647 4123 3684
rect 2414 2635 4122 2672
<< metal1 >>
rect 2418 3690 4121 3693
rect 2403 3684 4135 3690
rect 2403 3647 2415 3684
rect 4123 3647 4135 3684
rect 2403 3641 4135 3647
rect 2418 3625 4121 3641
rect 2790 3563 2834 3625
rect 2775 3510 2839 3563
rect 2971 3423 3010 3625
rect 3096 3514 3160 3567
rect 3407 3511 3471 3564
rect 2971 3384 3080 3423
rect 3146 3374 3250 3432
rect 2776 3282 2840 3335
rect 3094 3286 3158 3339
rect 3212 2934 3250 3374
rect 3182 2919 3250 2934
rect 3148 2918 3250 2919
rect 2960 2841 3027 2886
rect 1996 2618 2006 2700
rect 2080 2618 2090 2700
rect 2678 2693 2713 2794
rect 2960 2693 3005 2841
rect 3136 2832 3146 2918
rect 3204 2844 3250 2918
rect 3307 3393 3410 3432
rect 3542 3430 3581 3625
rect 3737 3566 3775 3625
rect 3728 3513 3792 3566
rect 3737 3509 3775 3513
rect 3307 2897 3346 3393
rect 3494 3391 3581 3430
rect 3408 3282 3472 3335
rect 3725 3284 3789 3337
rect 3307 2844 3319 2897
rect 3204 2832 3222 2844
rect 3148 2830 3222 2832
rect 3309 2830 3319 2844
rect 3392 2883 3402 2897
rect 3392 2844 3414 2883
rect 3546 2844 3601 2888
rect 3392 2830 3402 2844
rect 3062 2760 3516 2797
rect 3557 2693 3601 2844
rect 3834 2693 3864 2799
rect 2418 2678 4121 2693
rect 2402 2672 4134 2678
rect 2402 2635 2414 2672
rect 4122 2635 4134 2672
rect 2402 2629 4134 2635
rect 2418 2625 4121 2629
rect 5504 2372 5514 2448
rect 5598 2372 5608 2448
<< via1 >>
rect 2006 2618 2080 2700
rect 3146 2832 3204 2918
rect 3319 2830 3392 2897
rect 5514 2372 5598 2448
<< metal2 >>
rect 3146 2918 3204 2928
rect 3319 2897 3392 2907
rect 3146 2822 3204 2832
rect 3307 2830 3319 2857
rect 1986 2724 2100 2734
rect 3158 2678 3198 2822
rect 2100 2638 3198 2678
rect 3307 2820 3392 2830
rect 1986 2602 2100 2612
rect 3307 2614 3348 2820
rect 3307 2573 5598 2614
rect 5557 2468 5598 2573
rect 5484 2458 5600 2468
rect 5484 2346 5600 2356
<< via2 >>
rect 1986 2700 2100 2724
rect 1986 2618 2006 2700
rect 2006 2618 2080 2700
rect 2080 2618 2100 2700
rect 1986 2612 2100 2618
rect 5484 2448 5600 2458
rect 5484 2372 5514 2448
rect 5514 2372 5598 2448
rect 5598 2372 5600 2448
rect 5484 2356 5600 2372
<< metal3 >>
rect 1960 2608 1970 2748
rect 2120 2608 2130 2748
rect 1976 2607 2110 2608
rect 5474 2458 5610 2463
rect 5474 2356 5484 2458
rect 5600 2356 5610 2458
rect 5474 2351 5610 2356
<< via3 >>
rect 1970 2724 2120 2748
rect 1970 2612 1986 2724
rect 1986 2612 2100 2724
rect 2100 2612 2120 2724
rect 1970 2608 2120 2612
<< metal4 >>
rect 1969 2748 2121 2749
rect 1969 2608 1970 2748
rect 2120 2608 2121 2748
rect 1969 2607 2121 2608
rect 1994 2294 2054 2607
use sky130_fd_pr__cap_mim_m3_1_TNHPNJ  XC3
timestamp 1697379271
transform 1 0 3433 0 1 1481
box -2186 -1040 2186 1040
use sky130_fd_pr__nfet_01v8_SMGLWN  XM1
timestamp 1697915631
transform 1 0 3096 0 1 2881
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM2
timestamp 1697915631
transform 1 0 3482 0 1 2881
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_XJ7GBL  XM3
timestamp 1697379271
transform 1 0 3447 0 1 3424
box -211 -269 211 269
use sky130_fd_pr__nfet_01v8_SMGLWN  XM4
timestamp 1697915631
transform 1 0 2710 0 1 2881
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM5
timestamp 1697915631
transform 1 0 3868 0 1 2881
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_XJ7GBL  XM6
timestamp 1697379271
transform 1 0 2815 0 1 3424
box -211 -269 211 269
use sky130_fd_pr__pfet_01v8_XJ7GBL  XM7
timestamp 1697379271
transform 1 0 3763 0 1 3424
box -211 -269 211 269
use sky130_fd_pr__pfet_01v8_XJ7GBL  XM18
timestamp 1697379271
transform 1 0 3131 0 1 3424
box -211 -269 211 269
<< labels >>
rlabel metal2 4602 2614 4602 2614 1 vo1
rlabel metal1 4056 3693 4056 3693 1 Vdd
rlabel metal1 4134 2653 4134 2653 3 gnd
<< end >>
