magic
tech sky130A
magscale 1 2
timestamp 1699103691
<< dnwell >>
rect 124 38 1480 52
rect 124 -38 1738 38
rect 118 -1078 1738 -38
rect 124 -1092 1738 -1078
rect 124 -1118 1480 -1092
<< nwell >>
rect 1654 180 1896 182
rect -44 106 1896 180
rect -46 -68 1896 106
rect -46 -1012 242 -68
rect 498 -70 1896 -68
rect 1556 -1004 1896 -70
rect 1424 -1012 1896 -1004
rect -46 -1194 1896 -1012
rect -46 -1196 1672 -1194
rect 12 -1198 260 -1196
rect 1424 -1200 1672 -1196
<< nmos >>
rect 410 -766 610 -164
rect 1028 -762 1228 -160
<< ndiff >>
rect 350 -176 410 -164
rect 350 -752 364 -176
rect 398 -752 410 -176
rect 350 -764 410 -752
rect 352 -766 410 -764
rect 610 -176 668 -164
rect 610 -752 622 -176
rect 656 -752 668 -176
rect 610 -766 668 -752
rect 970 -174 1028 -160
rect 970 -750 982 -174
rect 1016 -750 1028 -174
rect 970 -762 1028 -750
rect 1228 -162 1286 -160
rect 1228 -174 1294 -162
rect 1228 -750 1240 -174
rect 1274 -750 1294 -174
rect 1228 -762 1294 -750
<< ndiffc >>
rect 364 -752 398 -176
rect 622 -752 656 -176
rect 982 -750 1016 -174
rect 1240 -750 1274 -174
<< psubdiff >>
rect 1390 -524 1512 -476
rect 1390 -786 1416 -524
rect 1476 -786 1512 -524
rect 1390 -860 1512 -786
<< nsubdiff >>
rect 1632 -530 1754 -470
rect 1632 -792 1656 -530
rect 1716 -792 1754 -530
rect 1632 -854 1754 -792
<< psubdiffcont >>
rect 1416 -786 1476 -524
<< nsubdiffcont >>
rect 1656 -792 1716 -530
<< poly >>
rect 410 -164 610 -136
rect 1028 -160 1228 -134
rect 410 -824 610 -766
rect 1028 -822 1228 -762
rect 1020 -824 1228 -822
rect 410 -840 630 -824
rect 410 -876 442 -840
rect 608 -876 630 -840
rect 410 -892 630 -876
rect 1008 -840 1228 -824
rect 1008 -874 1026 -840
rect 1186 -874 1228 -840
rect 1008 -892 1228 -874
<< polycont >>
rect 442 -876 608 -840
rect 1026 -874 1186 -840
<< locali >>
rect 346 -176 406 -158
rect 346 -752 364 -176
rect 398 -752 406 -176
rect 346 -768 406 -752
rect 606 -176 672 -154
rect 606 -752 622 -176
rect 656 -752 672 -176
rect 606 -770 672 -752
rect 982 -174 1016 -158
rect 982 -766 1016 -750
rect 1240 -174 1280 -158
rect 1274 -750 1280 -174
rect 1392 -476 1752 -472
rect 1240 -766 1280 -750
rect 1390 -524 1752 -476
rect 1390 -786 1416 -524
rect 1476 -530 1752 -524
rect 1476 -786 1656 -530
rect 1390 -792 1656 -786
rect 1716 -792 1752 -530
rect 1020 -824 1228 -822
rect 410 -840 630 -824
rect 410 -876 442 -840
rect 608 -876 630 -840
rect 410 -892 630 -876
rect 1008 -840 1228 -824
rect 1008 -874 1026 -840
rect 1186 -874 1228 -840
rect 1390 -856 1752 -792
rect 1390 -860 1512 -856
rect 1008 -892 1228 -874
<< viali >>
rect 364 -752 398 -176
rect 622 -752 656 -176
rect 982 -750 1016 -174
rect 1240 -750 1274 -174
rect 442 -876 608 -840
rect 1026 -874 1186 -840
<< metal1 >>
rect 346 -176 406 -158
rect 346 -752 364 -176
rect 398 -752 406 -176
rect 346 -768 406 -752
rect 606 -176 672 -154
rect 606 -752 622 -176
rect 656 -752 672 -176
rect 364 -935 398 -768
rect 606 -770 672 -752
rect 976 -174 1024 -162
rect 976 -750 982 -174
rect 1016 -750 1024 -174
rect 976 -762 1024 -750
rect 1234 -174 1282 -162
rect 1234 -750 1240 -174
rect 1274 -750 1282 -174
rect 1234 -762 1282 -750
rect 622 -824 656 -770
rect 982 -824 1016 -762
rect 1239 -766 1277 -762
rect 426 -840 656 -824
rect 426 -876 442 -840
rect 608 -876 656 -840
rect 426 -892 656 -876
rect 978 -840 1208 -824
rect 978 -874 1026 -840
rect 1186 -874 1208 -840
rect 978 -892 1208 -874
rect 1239 -884 1273 -766
rect 1239 -934 1272 -884
rect 756 -935 898 -934
rect 1238 -935 1272 -934
rect 364 -969 1272 -935
rect 364 -972 440 -969
rect 1238 -970 1272 -969
<< end >>
