magic
tech sky130A
magscale 1 2
timestamp 1699130246
<< nwell >>
rect 25622 1886 25868 2196
rect 7840 300 8660 626
rect 24460 464 24478 776
rect 15742 188 16140 428
rect 17918 192 18198 430
rect 19090 196 19372 430
rect 19948 428 24478 464
rect 19948 186 24476 428
<< poly >>
rect 1446 6970 1566 7098
rect 1412 6940 1566 6970
rect 1446 6778 1566 6940
rect 1414 6770 1566 6778
rect 1414 6748 1704 6770
rect 1444 6586 1704 6748
rect 1414 6556 1704 6586
rect 1444 6394 1704 6556
rect 1414 6364 1704 6394
rect 1444 6202 1704 6364
rect 1414 6172 1704 6202
rect 1444 6010 1704 6172
rect 1416 5980 1704 6010
rect 1444 5818 1704 5980
rect 1414 5788 1704 5818
rect 1444 5626 1704 5788
rect 1416 5596 1704 5626
rect 1444 5418 1704 5596
rect 1412 5388 1704 5418
rect 1444 5226 1704 5388
rect 1416 5196 1704 5226
rect 1444 5034 1704 5196
rect 1414 5004 1704 5034
rect 1444 4938 1704 5004
rect 1410 4908 1704 4938
rect 1444 4842 1704 4908
rect 1408 4812 1704 4842
rect 1444 4650 1704 4812
rect 1410 4620 1704 4650
rect 1444 4458 1704 4620
rect 1408 4428 1704 4458
rect 1444 4266 1704 4428
rect 1414 4236 1704 4266
rect 1444 4074 1704 4236
rect 1408 4044 1704 4074
rect 1444 3882 1704 4044
rect 1408 3852 1704 3882
rect 1444 3690 1704 3852
rect 1408 3660 1704 3690
rect 1444 3498 1704 3660
rect 1410 3468 1704 3498
rect 1444 3306 1704 3468
rect 1408 3276 1704 3306
rect 1444 3114 1704 3276
rect 1408 3084 1704 3114
rect 1444 2922 1704 3084
rect 1408 2892 1704 2922
rect 1444 2730 1704 2892
rect 1406 2700 1704 2730
rect 1444 2538 1704 2700
rect 1408 2508 1704 2538
rect 1444 2346 1704 2508
rect 1408 2316 1704 2346
rect 1444 2154 1704 2316
rect 1408 2124 1704 2154
rect 1444 1962 1704 2124
rect 1410 1932 1704 1962
rect 1444 1770 1704 1932
rect 1410 1740 1704 1770
rect 1444 1578 1704 1740
rect 1408 1548 1704 1578
rect 1444 1386 1704 1548
rect 1408 1356 1704 1386
rect 1444 1194 1704 1356
rect 1410 1164 1704 1194
rect 1444 1002 1704 1164
rect 1404 972 1704 1002
rect 1444 810 1704 972
rect 1412 780 1704 810
rect 1444 614 1704 780
rect 15768 326 16000 424
rect 17918 192 18198 430
<< locali >>
rect 1446 6838 1704 7098
rect 1444 6794 1704 6838
rect 1444 6708 1834 6794
rect 1444 742 1538 6708
rect 1730 742 1834 6708
rect 1444 614 1834 742
rect 15768 364 16000 424
rect 15738 326 16000 364
rect 15738 184 15994 326
rect 17918 192 18198 430
<< viali >>
rect 1538 742 1730 6708
<< metal1 >>
rect 1024 8002 1388 9242
rect 924 7938 1388 8002
rect 924 7584 990 7938
rect 1314 7584 1388 7938
rect 25308 8238 25734 8428
rect 924 7520 1388 7584
rect 1024 542 1388 7520
rect 1494 7366 1844 7676
rect 24596 7490 25130 7686
rect 1484 7320 2060 7366
rect 1484 7180 1514 7320
rect 2012 7180 2060 7320
rect 1484 7156 2060 7180
rect 24560 7344 25152 7490
rect 1494 6708 1844 7156
rect 24560 6930 24614 7344
rect 25062 6930 25152 7344
rect 25308 7288 25400 8238
rect 25612 7288 25734 8238
rect 25308 7000 25734 7288
rect 25622 6990 25734 7000
rect 24560 6866 25152 6930
rect 24596 6852 24722 6866
rect 1494 742 1538 6708
rect 1730 786 1844 6708
rect 23384 1092 23856 1094
rect 9546 1066 13142 1072
rect 7450 994 9094 1046
rect 7450 808 7532 994
rect 8980 808 9094 994
rect 1730 742 2598 786
rect 1494 612 2598 742
rect 7450 621 9094 808
rect 9380 1022 13142 1066
rect 9380 684 9422 1022
rect 9810 684 13142 1022
rect 9380 654 13142 684
rect 23384 1048 23872 1092
rect 23384 870 23440 1048
rect 23822 870 23872 1048
rect 9380 650 9860 654
rect 1494 604 1844 612
rect 7450 600 7991 621
rect 8208 600 9094 621
rect 8551 579 8591 600
rect 23384 590 23872 870
rect 23400 588 23872 590
rect 782 534 1408 542
rect 782 -40 6076 534
rect 9154 386 9514 422
rect 9154 252 9188 386
rect 7772 199 8520 232
rect 9016 219 9188 252
rect 7460 24 7494 86
rect 7678 32 7712 86
rect 7620 24 7714 32
rect 7460 21 7714 24
rect 7426 17 7714 21
rect 932 -470 6076 -40
rect 7456 4 7714 17
rect 7456 -10 8156 4
rect 8706 -10 8740 102
rect 8924 -10 8958 102
rect 9154 88 9188 219
rect 9462 88 9514 386
rect 9154 56 9514 88
rect 7456 -56 8966 -10
rect 7456 -262 7522 -56
rect 8864 -262 8966 -56
rect 7456 -302 8966 -262
rect 9632 -110 13100 524
rect 17918 428 18198 430
rect 15742 188 16140 428
rect 17838 200 18326 428
rect 17918 192 18198 200
rect 9632 -422 9690 -110
rect 10684 -422 13100 -110
rect 24320 -102 24914 384
rect 24320 -364 24382 -102
rect 24834 -364 24914 -102
rect 24320 -412 24914 -364
rect 9632 -462 13100 -422
rect 9636 -464 10774 -462
<< via1 >>
rect 990 7584 1314 7938
rect 1514 7180 2012 7320
rect 24614 6930 25062 7344
rect 25400 7288 25612 8238
rect 7532 808 8980 994
rect 9422 684 9810 1022
rect 23440 870 23822 1048
rect 9188 88 9462 386
rect 7522 -262 8864 -56
rect 9690 -422 10684 -110
rect 24382 -364 24834 -102
<< metal2 >>
rect 25316 8238 25682 8354
rect 924 7938 1368 8002
rect 924 7584 990 7938
rect 1314 7584 1368 7938
rect 924 7520 1368 7584
rect 24560 7490 25132 7494
rect 1484 7320 2060 7366
rect 1484 7180 1514 7320
rect 2012 7180 2060 7320
rect 1484 7156 2060 7180
rect 24560 7344 25152 7490
rect 24560 6930 24614 7344
rect 25062 6930 25152 7344
rect 25316 7288 25400 8238
rect 25612 7288 25682 8238
rect 25316 7246 25682 7288
rect 24560 6866 25152 6930
rect 24560 6862 24722 6866
rect 7458 1046 7818 1048
rect 7458 994 9078 1046
rect 7458 808 7532 994
rect 8980 808 9078 994
rect 7458 756 9078 808
rect 9380 1022 9860 1066
rect 7458 748 7818 756
rect 9380 684 9422 1022
rect 9810 684 9860 1022
rect 23380 1048 23894 1096
rect 23380 870 23440 1048
rect 23822 870 23894 1048
rect 23380 798 23894 870
rect 9380 650 9860 684
rect 6586 402 7258 426
rect 6586 78 6648 402
rect 7052 317 7258 402
rect 9154 386 9514 422
rect 7052 111 7391 317
rect 7052 78 7258 111
rect 6586 52 7258 78
rect 9154 88 9188 386
rect 9462 88 9514 386
rect 9154 56 9514 88
rect 7456 -56 8966 -10
rect 7456 -262 7522 -56
rect 8864 -262 8966 -56
rect 7456 -302 8966 -262
rect 9636 -110 10774 -58
rect 9636 -422 9690 -110
rect 10684 -422 10774 -110
rect 24320 -102 24918 -30
rect 24320 -364 24382 -102
rect 24834 -364 24918 -102
rect 24320 -412 24918 -364
rect 9636 -464 10774 -422
<< via2 >>
rect 990 7584 1314 7938
rect 1514 7180 2012 7320
rect 24614 6930 25062 7344
rect 25400 7288 25612 8238
rect 7532 808 8980 994
rect 9422 684 9810 1022
rect 23440 870 23822 1048
rect 6648 78 7052 402
rect 9188 88 9462 386
rect 7522 -262 8864 -56
rect 9690 -422 10684 -110
rect 24382 -364 24834 -102
<< metal3 >>
rect 25316 8238 25682 8354
rect 924 7938 1368 8002
rect 924 7584 990 7938
rect 1314 7584 1368 7938
rect 924 7520 1368 7584
rect 24560 7490 25132 7494
rect 1484 7320 2060 7366
rect 1484 7180 1514 7320
rect 2012 7180 2060 7320
rect 1484 7156 2060 7180
rect 24560 7344 25152 7490
rect 24560 6930 24614 7344
rect 25062 6930 25152 7344
rect 25316 7288 25400 8238
rect 25612 7288 25682 8238
rect 25316 7246 25682 7288
rect 24560 6866 25152 6930
rect 24560 6862 24722 6866
rect 7458 1046 7818 1048
rect 7458 994 9078 1046
rect 7458 808 7532 994
rect 8980 808 9078 994
rect 7458 756 9078 808
rect 9380 1022 9860 1066
rect 7458 748 7818 756
rect 9380 684 9422 1022
rect 9810 684 9860 1022
rect 9380 650 9860 684
rect 6586 424 7258 426
rect 13297 424 13431 2597
rect 23380 1048 23894 1096
rect 23380 870 23440 1048
rect 23822 870 23894 1048
rect 23380 798 23894 870
rect 1805 402 7258 424
rect 1805 78 6648 402
rect 7052 78 7258 402
rect 1805 52 7258 78
rect 9144 386 25666 424
rect 9144 88 9188 386
rect 9462 332 25666 386
rect 9462 88 25447 332
rect 1805 46 6916 52
rect 9144 46 25447 88
rect 7456 -56 8966 -10
rect 7456 -262 7522 -56
rect 8864 -262 8966 -56
rect 7456 -302 8966 -262
rect 9636 -110 10774 -58
rect 9636 -422 9690 -110
rect 10684 -422 10774 -110
rect 24320 -102 24918 -30
rect 24320 -364 24382 -102
rect 24834 -364 24918 -102
rect 24320 -412 24918 -364
rect 9636 -464 10774 -422
<< via3 >>
rect 990 7584 1314 7938
rect 1514 7180 2012 7320
rect 24614 6930 25062 7344
rect 25400 7288 25612 8238
rect 7532 808 8980 994
rect 9422 684 9810 1022
rect 23440 870 23822 1048
rect 7522 -262 8864 -56
rect 9690 -422 10684 -110
rect 24382 -364 24834 -102
<< metal4 >>
rect 25316 8266 25682 8354
rect 924 7938 1368 8002
rect 924 7584 990 7938
rect 1314 7584 1368 7938
rect 924 7520 1368 7584
rect 1484 7320 2060 7366
rect 1484 7180 1514 7320
rect 2012 7180 2060 7320
rect 1484 7156 2060 7180
rect 24560 7344 25160 7494
rect 24560 7086 24614 7344
rect 24554 6930 24614 7086
rect 25062 6930 25160 7344
rect 25316 7288 25400 8266
rect 25640 8230 25682 8266
rect 25648 7288 25682 8230
rect 25316 7246 25682 7288
rect 1488 1136 2056 5158
rect 24554 1136 25160 6930
rect 1488 1048 25160 1136
rect 1488 1022 23440 1048
rect 1488 994 9422 1022
rect 1488 808 7532 994
rect 8980 808 9422 994
rect 1488 684 9422 808
rect 9810 870 23440 1022
rect 23822 870 25160 1048
rect 9810 684 25160 870
rect 1488 578 25160 684
rect 1488 568 24670 578
rect 7456 -28 8966 -10
rect 7456 -276 7518 -28
rect 8874 -276 8966 -28
rect 7456 -302 8966 -276
rect 9636 -110 10774 -58
rect 9636 -422 9690 -110
rect 10684 -422 10774 -110
rect 24320 -102 24918 -30
rect 24320 -364 24382 -102
rect 24834 -364 24918 -102
rect 24320 -412 24918 -364
rect 9636 -464 10774 -422
<< via4 >>
rect 990 7584 1314 7938
rect 25400 8238 25640 8266
rect 25400 7288 25612 8238
rect 25612 8230 25640 8238
rect 25612 7288 25648 8230
rect 7518 -56 8874 -28
rect 7518 -262 7522 -56
rect 7522 -262 8864 -56
rect 8864 -262 8874 -56
rect 7518 -276 8874 -262
rect 9690 -422 10684 -110
rect 24382 -364 24834 -102
<< metal5 >>
rect 789 7938 1393 10802
rect 789 7584 990 7938
rect 1314 7584 1393 7938
rect 789 46 1393 7584
rect 25314 7288 25400 7877
rect 25648 7288 25904 7877
rect 25314 46 25904 7288
rect 789 -28 25904 46
rect 789 -276 7518 -28
rect 8874 -102 25904 -28
rect 8874 -110 24382 -102
rect 8874 -276 9690 -110
rect 789 -422 9690 -276
rect 10684 -364 24382 -110
rect 24834 -364 25904 -102
rect 10684 -422 25904 -364
rect 789 -507 25904 -422
rect 789 -558 25892 -507
use buffer_digital  buffer_digital_0
timestamp 1699114361
transform 1 0 8708 0 1 68
box -274 -35 412 578
use buffer_digital  buffer_digital_1
timestamp 1699114361
transform 1 0 7462 0 1 52
box -274 -35 412 578
use charge_pump1  charge_pump1_0
timestamp 1699130246
transform 1 0 821 0 1 10004
box -313 -7588 25321 19132
use nmos_decap_10  nmos_decap_10_0
timestamp 1699103691
transform 1 0 2110 0 1 368
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_1
timestamp 1699103691
transform 1 0 3070 0 1 368
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_2
timestamp 1699103691
transform 1 0 4030 0 1 368
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_3
timestamp 1699103691
transform 1 0 4990 0 1 368
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_4
timestamp 1699103691
transform 1 0 10022 0 1 366
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_5
timestamp 1699103691
transform 1 0 10982 0 1 366
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_6
timestamp 1699103691
transform 1 0 11942 0 1 366
box -10 -42 1060 416
use pmos_decap_10  pmos_decap_10_0
timestamp 1699103691
transform 1 0 13704 0 -1 650
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_1
timestamp 1699103691
transform -1 0 15874 0 -1 652
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_2
timestamp 1699103691
transform 1 0 15862 0 -1 654
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_3
timestamp 1699103691
transform -1 0 18034 0 -1 658
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_4
timestamp 1699103691
transform 1 0 18016 0 -1 658
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_5
timestamp 1699103691
transform 1 0 19090 0 -1 660
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_6
timestamp 1699103691
transform 1 0 20162 0 -1 670
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_7
timestamp 1699103691
transform 1 0 21234 0 -1 666
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_8
timestamp 1699103691
transform 1 0 22306 0 -1 666
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_9
timestamp 1699103691
transform 1 0 23380 0 -1 670
box 0 -108 1098 464
use sky130_fd_pr__nfet_01v8_HRDN5X  sky130_fd_pr__nfet_01v8_HRDN5X_0
timestamp 1699103691
transform 0 1 1364 -1 0 6283
box -749 -130 749 130
use sky130_fd_pr__nfet_01v8_TKGCLY  sky130_fd_pr__nfet_01v8_TKGCLY_0
timestamp 1699103691
transform 0 1 1358 -1 0 3051
box -2429 -130 2429 130
<< labels >>
rlabel metal3 6365 145 6365 145 1 clk_in
rlabel metal3 9567 169 9567 169 1 clk_out
rlabel metal1 8130 206 8130 206 1 clk_int
rlabel metal4 7299 650 7299 650 1 vdd
rlabel metal5 7313 -49 7313 -49 1 gnd
<< end >>
