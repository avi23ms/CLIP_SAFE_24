magic
tech sky130A
magscale 1 2
timestamp 1698179620
<< pwell >>
rect 610 3878 694 3892
rect -2830 3732 -2512 3810
rect 126 3732 406 3842
rect 608 3738 694 3878
rect 610 3724 694 3738
rect 3440 3726 3880 3840
rect -1219 3461 -1134 3531
<< locali >>
rect 488 4848 562 4932
rect 474 3738 562 3830
rect 474 3730 600 3738
rect -849 3234 -790 3381
rect -2215 2557 -1907 2591
rect -1827 2545 -1682 2579
rect -1440 2562 -1295 2596
rect -1059 2549 -751 2583
rect -2032 2386 -1991 2491
rect -867 2386 -826 2491
rect -2255 2365 -599 2386
rect -2255 2308 -599 2325
<< viali >>
rect -2255 2325 -599 2365
<< metal1 >>
rect -2922 5468 -2720 5522
rect 3792 5468 3966 5482
rect -3704 5304 -3694 5468
rect 4116 5304 4126 5468
rect -2922 5178 -2720 5304
rect -2918 4918 -2720 5178
rect -3163 4836 -2720 4918
rect -3163 3495 -3081 4836
rect -2918 4791 -2720 4836
rect 3792 4826 3966 5304
rect 54 4678 64 4744
rect 152 4678 162 4744
rect 3506 4678 3516 4738
rect 3622 4678 3632 4738
rect -1190 4552 -1180 4632
rect -1102 4552 -1092 4632
rect -3042 3945 -2810 3986
rect -3042 3580 -3001 3945
rect -2766 3736 -2756 3790
rect -2524 3736 -2514 3790
rect -1921 3666 -1817 3684
rect -1922 3604 -1912 3666
rect -1836 3664 -1817 3666
rect -1921 3585 -1890 3604
rect -3042 3539 -1955 3580
rect -3163 3413 -2225 3495
rect -2307 2386 -2225 3413
rect -1996 2904 -1955 3539
rect -1914 2970 -1890 3585
rect -1834 3585 -1817 3664
rect -1352 3620 -1302 3766
rect 118 3734 128 3786
rect 380 3734 390 3786
rect 602 3718 612 3792
rect 688 3718 698 3792
rect 3436 3724 3446 3808
rect 3778 3724 3788 3808
rect -1834 2998 -1818 3585
rect -1185 3575 -1147 3595
rect -1185 3535 -945 3575
rect -655 3570 -620 3614
rect -1253 3529 -945 3535
rect -1253 3497 -1134 3529
rect -670 3528 1508 3570
rect -1426 3461 -1134 3497
rect -655 3476 -586 3528
rect -1426 3460 -1135 3461
rect -1253 3457 -1135 3460
rect -655 3129 -618 3476
rect 3674 3262 3684 3264
rect 3364 3200 3400 3262
rect 3480 3200 3546 3262
rect 3626 3202 3684 3262
rect 3764 3262 3774 3264
rect 3764 3260 3888 3262
rect 3764 3202 3802 3260
rect 3626 3200 3802 3202
rect 3792 3198 3802 3200
rect 3882 3198 3892 3260
rect -1251 3061 -697 3098
rect -1834 2990 -1112 2998
rect -1834 2970 1286 2990
rect -1914 2961 1286 2970
rect -1149 2958 1286 2961
rect -2006 2830 -1996 2904
rect -1551 2822 -1541 2830
rect -1452 2822 -1442 2904
rect -1712 2672 -1702 2740
rect -1594 2672 -1584 2740
rect -1542 2544 -1501 2822
rect -1149 2542 -1112 2958
rect -630 2802 -620 2892
rect -530 2802 -520 2892
rect -462 2816 -452 2878
rect -390 2816 -380 2878
rect -312 2822 -302 2884
rect -240 2822 -230 2884
rect -180 2822 -170 2884
rect -108 2822 -98 2884
rect -46 2822 -36 2884
rect 26 2822 36 2884
rect 1254 2662 1286 2958
rect 1254 2630 1874 2662
rect 1842 2532 1874 2630
rect 2162 2530 2172 2584
rect 2238 2530 2248 2584
rect -1683 2433 -1673 2495
rect -1566 2481 -1556 2495
rect -1566 2452 -1201 2481
rect -1566 2433 -1556 2452
rect -2307 2381 -599 2386
rect -2307 2365 -131 2381
rect -2307 2325 -2255 2365
rect -599 2325 -131 2365
rect -2432 2259 -2422 2320
rect -2362 2259 -2352 2320
rect -2307 2299 -131 2325
rect -213 1883 -131 2299
rect 402 2166 412 2318
rect 570 2166 580 2318
rect 694 2168 704 2314
rect 854 2168 864 2314
rect 4250 2208 4680 2256
rect -213 1824 -193 1883
rect -130 1824 -120 1883
rect -213 1716 -131 1824
rect 4276 1770 4286 1840
rect 4354 1770 4364 1840
rect -213 1660 -188 1716
rect -128 1660 -118 1716
rect -213 1608 -131 1660
rect 4278 1614 4288 1700
rect 4354 1614 4364 1700
rect -213 1552 -190 1608
rect -130 1552 -120 1608
rect -213 1478 -131 1552
rect -213 1422 -190 1478
rect -130 1422 -120 1478
rect 4278 1456 4288 1542
rect 4354 1456 4364 1542
rect -213 1352 -131 1422
rect -213 1296 -188 1352
rect -128 1296 -118 1352
rect -213 1206 -131 1296
rect 4274 1282 4284 1368
rect 4350 1282 4360 1368
rect -213 1150 -188 1206
rect -128 1150 -118 1206
rect -213 77 -131 1150
rect 4278 1094 4288 1180
rect 4354 1094 4364 1180
rect 4632 -176 4680 2208
rect -3568 -404 4956 -176
rect -3578 -654 -3568 -404
rect 4922 -654 4956 -404
rect -3568 -810 4956 -654
<< via1 >>
rect -3694 5304 4116 5468
rect 64 4678 152 4744
rect 3516 4678 3622 4738
rect -1180 4552 -1102 4632
rect -2756 3736 -2524 3790
rect -1912 3664 -1836 3666
rect -1912 3604 -1834 3664
rect -1890 2970 -1834 3604
rect 128 3734 380 3786
rect 612 3718 688 3792
rect 3446 3724 3778 3808
rect 3400 3200 3480 3262
rect 3546 3200 3626 3262
rect 3684 3202 3764 3264
rect 3802 3198 3882 3260
rect -1996 2830 -1452 2904
rect -1541 2822 -1452 2830
rect -1702 2672 -1594 2740
rect -620 2802 -530 2892
rect -452 2816 -390 2878
rect -302 2822 -240 2884
rect -170 2822 -108 2884
rect -36 2822 26 2884
rect 2172 2530 2238 2584
rect -1673 2433 -1566 2495
rect -2422 2259 -2362 2320
rect 412 2166 570 2318
rect 704 2168 854 2314
rect -193 1824 -130 1883
rect 4286 1770 4354 1840
rect -188 1660 -128 1716
rect 4288 1614 4354 1700
rect -190 1552 -130 1608
rect -190 1422 -130 1478
rect 4288 1456 4354 1542
rect -188 1296 -128 1352
rect 4284 1282 4350 1368
rect -188 1150 -128 1206
rect 4288 1094 4354 1180
rect -3568 -654 4922 -404
<< metal2 >>
rect -3694 5468 4116 5478
rect -3694 5294 4116 5304
rect -3283 5005 -1134 5043
rect -3283 2764 -3245 5005
rect -1172 4642 -1134 5005
rect 68 4998 3572 5054
rect 68 4754 124 4998
rect 64 4744 152 4754
rect 64 4668 152 4678
rect 3516 4748 3572 4998
rect 3516 4738 3622 4748
rect 3516 4668 3622 4678
rect -1180 4632 -1102 4642
rect -1180 4542 -1102 4552
rect -2828 3837 -2785 3915
rect -2828 3810 -2750 3837
rect -2830 3790 -2512 3810
rect -2830 3736 -2756 3790
rect -2524 3736 -2512 3790
rect -2830 3732 -2512 3736
rect -2756 3726 -2524 3732
rect -2189 3672 -2147 4199
rect 350 3842 392 3923
rect 610 3878 694 3892
rect 126 3786 406 3842
rect 126 3734 128 3786
rect 380 3734 406 3786
rect 608 3792 694 3878
rect 608 3738 612 3792
rect 126 3732 406 3734
rect 128 3724 380 3732
rect 610 3724 612 3738
rect 688 3724 694 3792
rect 612 3708 688 3718
rect -1912 3674 -1836 3676
rect -1912 3672 -1834 3674
rect -2192 3666 -1834 3672
rect -2192 3630 -1912 3666
rect -1836 3664 -1834 3666
rect -1912 3594 -1890 3604
rect -1890 2960 -1834 2970
rect -1996 2904 -1452 2914
rect -620 2892 -530 2902
rect -1996 2822 -1541 2830
rect -1452 2822 -620 2878
rect -1996 2820 -1452 2822
rect -1541 2812 -1452 2820
rect -452 2878 -390 2888
rect -302 2884 -240 2894
rect -530 2822 -452 2878
rect -390 2822 -302 2878
rect -170 2884 -108 2894
rect -240 2822 -170 2878
rect -36 2884 26 2894
rect -108 2822 -36 2878
rect 26 2822 112 2878
rect -452 2806 -390 2816
rect -302 2812 -240 2822
rect -170 2812 -108 2822
rect -36 2812 26 2822
rect -620 2792 -530 2802
rect -3283 2750 -1614 2764
rect -3283 2740 -1594 2750
rect -3283 2728 -1702 2740
rect -3283 2727 -3245 2728
rect -1702 2662 -1594 2672
rect -1673 2495 -1566 2505
rect -2367 2442 -1673 2481
rect -2367 2341 -2328 2442
rect -1673 2423 -1566 2433
rect 838 2394 918 3962
rect 3816 3840 3858 3937
rect 3440 3808 3880 3840
rect 3440 3726 3446 3808
rect 3778 3726 3880 3808
rect 3446 3714 3778 3724
rect 3400 3262 3480 3272
rect 3400 3190 3480 3200
rect 3546 3262 3626 3272
rect 3546 3190 3626 3200
rect 3684 3264 3764 3274
rect 3684 3192 3764 3202
rect 3802 3260 3882 3270
rect 3802 3188 3882 3198
rect 2172 2588 2238 2598
rect 2172 2520 2238 2530
rect -2442 2331 -2328 2341
rect -2340 2285 -2328 2331
rect 412 2318 570 2328
rect 798 2324 920 2394
rect -2442 2232 -2340 2242
rect 264 2168 412 2308
rect 264 2164 322 2168
rect 704 2314 920 2324
rect 570 2168 704 2308
rect 854 2308 920 2314
rect 854 2168 1146 2308
rect 412 2156 570 2166
rect 704 2158 854 2168
rect -213 1890 -129 1900
rect 4310 1850 4351 2164
rect -213 1796 -129 1806
rect 4286 1840 4354 1850
rect 4286 1760 4354 1770
rect -188 1716 -128 1726
rect 4310 1710 4351 1760
rect -188 1650 -128 1660
rect 4288 1700 4354 1710
rect -190 1608 -130 1618
rect 4288 1604 4354 1614
rect 4310 1552 4351 1604
rect -190 1542 -130 1552
rect 4288 1542 4354 1552
rect -190 1478 -130 1488
rect 4288 1446 4354 1456
rect -190 1412 -130 1422
rect 4310 1378 4351 1446
rect 4284 1368 4351 1378
rect -188 1352 -128 1362
rect -188 1286 -128 1296
rect 4350 1282 4351 1368
rect 4284 1272 4351 1282
rect -188 1206 -128 1216
rect 4310 1190 4351 1272
rect -188 1140 -128 1150
rect 4288 1180 4354 1190
rect 4288 1084 4354 1094
rect 4310 18 4351 1084
rect -3568 -404 4922 -394
rect -3568 -664 4922 -654
<< via2 >>
rect -3694 5304 4116 5468
rect -620 2802 -530 2892
rect -452 2816 -390 2878
rect -302 2822 -240 2884
rect -170 2822 -108 2884
rect -36 2822 26 2884
rect 2172 2584 2238 2588
rect 2172 2530 2238 2584
rect -2442 2320 -2340 2331
rect -2442 2259 -2422 2320
rect -2422 2259 -2362 2320
rect -2362 2259 -2340 2320
rect -2442 2242 -2340 2259
rect 412 2166 570 2318
rect 704 2168 854 2314
rect -213 1883 -129 1890
rect -213 1824 -193 1883
rect -193 1824 -130 1883
rect -130 1824 -129 1883
rect -213 1806 -129 1824
rect 4286 1770 4354 1840
rect -188 1660 -128 1716
rect -190 1552 -130 1608
rect 4288 1614 4354 1700
rect -190 1422 -130 1478
rect 4288 1456 4354 1542
rect -188 1296 -128 1352
rect 4284 1282 4350 1368
rect -188 1150 -128 1206
rect 4288 1094 4354 1180
rect -3568 -654 4922 -404
<< metal3 >>
rect -3704 5304 -3694 5520
rect 4100 5473 4110 5520
rect 4100 5468 4126 5473
rect 4116 5304 4126 5468
rect -3704 5299 4126 5304
rect -538 2897 -470 2900
rect -630 2896 -470 2897
rect -630 2892 2262 2896
rect -630 2802 -620 2892
rect -530 2884 2262 2892
rect -530 2878 -302 2884
rect -530 2816 -452 2878
rect -390 2822 -302 2878
rect -240 2822 -170 2884
rect -108 2822 -36 2884
rect 26 2866 2262 2884
rect 26 2822 2266 2866
rect -390 2816 2266 2822
rect -530 2806 2266 2816
rect -530 2802 -470 2806
rect -630 2797 -470 2802
rect -538 2792 -470 2797
rect 2154 2588 2266 2806
rect 2154 2530 2172 2588
rect 2238 2530 2266 2588
rect 2162 2525 2248 2530
rect -2474 2214 -2464 2376
rect -2314 2214 -2304 2376
rect 402 2318 580 2323
rect 402 2310 412 2318
rect 136 2166 412 2310
rect 570 2310 580 2318
rect 694 2314 864 2319
rect 694 2310 704 2314
rect 570 2168 704 2310
rect 854 2310 864 2314
rect 854 2168 990 2310
rect 570 2166 990 2168
rect 402 2161 580 2166
rect 694 2163 864 2166
rect -223 1890 -119 1895
rect -223 1806 -213 1890
rect -129 1806 -119 1890
rect -223 1801 -119 1806
rect 4276 1840 4364 1845
rect 4276 1770 4286 1840
rect 4354 1770 4364 1840
rect 4276 1765 4364 1770
rect -198 1716 -118 1721
rect -198 1660 -188 1716
rect -128 1660 -118 1716
rect -198 1655 -118 1660
rect 4278 1700 4364 1705
rect 4278 1614 4288 1700
rect 4354 1614 4364 1700
rect -200 1608 -120 1613
rect 4278 1609 4364 1614
rect -200 1552 -190 1608
rect -130 1552 -120 1608
rect -200 1547 -120 1552
rect 4278 1542 4364 1547
rect -200 1478 -120 1483
rect -200 1422 -190 1478
rect -130 1422 -120 1478
rect 4278 1456 4288 1542
rect 4354 1456 4364 1542
rect 4278 1451 4364 1456
rect -200 1417 -120 1422
rect 4274 1368 4360 1373
rect -198 1352 -118 1357
rect -198 1296 -188 1352
rect -128 1296 -118 1352
rect -198 1291 -118 1296
rect 4274 1282 4284 1368
rect 4350 1282 4360 1368
rect 4274 1277 4360 1282
rect -198 1206 -118 1211
rect -198 1150 -188 1206
rect -128 1150 -118 1206
rect -198 1145 -118 1150
rect 4278 1180 4364 1185
rect 4278 1094 4288 1180
rect 4354 1094 4364 1180
rect 4278 1089 4364 1094
rect -3578 -654 -3568 -362
rect 4918 -399 4928 -362
rect 4918 -404 4932 -399
rect 4922 -654 4932 -404
rect -3578 -659 4932 -654
<< via3 >>
rect -3694 5468 4100 5520
rect -3694 5304 4100 5468
rect -2464 2331 -2314 2376
rect -2464 2242 -2442 2331
rect -2442 2242 -2340 2331
rect -2340 2242 -2314 2331
rect -2464 2214 -2314 2242
rect 412 2166 570 2318
rect 704 2168 854 2314
rect -3568 -404 4918 -362
rect -3568 -654 4922 -404
<< metal4 >>
rect -3694 5521 4108 5598
rect -3695 5520 4108 5521
rect -3695 5304 -3694 5520
rect 4100 5304 4108 5520
rect -3695 5303 4108 5304
rect -3694 5224 4108 5303
rect -2478 2376 -2296 2382
rect -2478 2214 -2464 2376
rect -2314 2214 -2296 2376
rect 411 2318 571 2319
rect 411 2312 412 2318
rect 136 2306 412 2312
rect -2478 1954 -2296 2214
rect 128 2166 412 2306
rect 570 2312 571 2318
rect 703 2314 855 2315
rect 703 2312 704 2314
rect 570 2168 704 2312
rect 854 2312 855 2314
rect 854 2168 1140 2312
rect 570 2166 1140 2168
rect -2478 1550 -2300 1954
rect 128 1902 292 2166
rect 411 2165 571 2166
rect -3569 -362 4919 -361
rect -3569 -654 -3568 -362
rect 4918 -403 4919 -362
rect 4918 -404 4923 -403
rect 4922 -654 4923 -404
rect -3569 -655 4923 -654
<< via4 >>
rect -3568 -654 4918 -362
<< metal5 >>
rect -3584 -338 4954 -174
rect -3592 -362 4954 -338
rect -3592 -654 -3568 -362
rect 4918 -654 4954 -362
rect -3592 -678 4954 -654
rect -3584 -808 4954 -678
use cmfb  cmfb_0
timestamp 1698179620
transform 1 0 -3134 0 1 2875
box 203 439 3639 2056
use integrator_full_new1  integrator_full_new1_0
timestamp 1698179620
transform 1 0 386 0 1 3314
box -386 -3314 3986 1624
use sky130_fd_pr__nfet_01v8_53744R  sky130_fd_pr__nfet_01v8_53744R_0
timestamp 1698166690
transform 0 1 -809 -1 0 3174
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_53744R  sky130_fd_pr__nfet_01v8_53744R_1
timestamp 1698166690
transform 0 1 -1323 -1 0 3560
box -246 -310 246 310
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_0
timestamp 1698155087
transform 1 0 -1233 0 1 2582
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_1
timestamp 1698155087
transform 1 0 -1619 0 1 2582
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_2
timestamp 1698155087
transform 1 0 -2005 0 1 2582
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_3
timestamp 1698155087
transform 1 0 -847 0 1 2582
box -246 -269 246 269
use sky130_fd_pr__cap_mim_m3_1_4PHTN9  XC3
timestamp 1697610037
transform 1 0 -1291 0 1 1094
box -1186 -1040 1186 1040
<< end >>
