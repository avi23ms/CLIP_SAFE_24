magic
tech sky130A
magscale 1 2
timestamp 1698837094
<< nwell >>
rect 7840 300 8660 626
<< nsubdiff >>
rect 8012 524 8190 548
rect 8012 370 8038 524
rect 8154 370 8190 524
rect 8012 352 8190 370
<< nsubdiffcont >>
rect 8038 370 8154 524
<< locali >>
rect 8012 524 8190 548
rect 8012 370 8038 524
rect 8154 370 8190 524
rect 8012 352 8190 370
<< viali >>
rect 8038 370 8154 524
<< metal1 >>
rect 7450 994 9094 1046
rect 7450 808 7532 994
rect 8980 808 9094 994
rect 7450 600 9094 808
rect 8036 548 8156 600
rect 8012 524 8190 548
rect 8012 370 8038 524
rect 8154 370 8190 524
rect 8012 352 8190 370
rect 9154 386 9514 422
rect 9154 252 9188 386
rect 7815 199 8520 232
rect 9016 219 9188 252
rect 7460 -10 7494 86
rect 7678 -10 7712 86
rect 8706 -10 8740 102
rect 8924 -10 8958 102
rect 9154 88 9188 219
rect 9462 88 9514 386
rect 9154 56 9514 88
rect 7456 -56 8966 -10
rect 7456 -262 7522 -56
rect 8864 -262 8966 -56
rect 7456 -302 8966 -262
<< via1 >>
rect 7532 808 8980 994
rect 9188 88 9462 386
rect 7522 -262 8864 -56
<< metal2 >>
rect 7458 1046 7818 1048
rect 7458 994 9078 1046
rect 7458 808 7532 994
rect 8980 808 9078 994
rect 7458 756 9078 808
rect 7458 748 7818 756
rect 6586 402 7258 426
rect 6586 78 6648 402
rect 7052 317 7258 402
rect 9154 386 9514 422
rect 7052 111 7391 317
rect 7052 78 7258 111
rect 6586 52 7258 78
rect 9154 88 9188 386
rect 9462 88 9514 386
rect 9154 56 9514 88
rect 7456 -56 8966 -10
rect 7456 -262 7522 -56
rect 8864 -262 8966 -56
rect 7456 -302 8966 -262
<< via2 >>
rect 7532 808 8980 994
rect 6648 78 7052 402
rect 9188 88 9462 386
rect 7522 -262 8864 -56
<< metal3 >>
rect 7458 1046 7818 1048
rect 7458 994 9078 1046
rect 7458 808 7532 994
rect 8980 808 9078 994
rect 7458 756 9078 808
rect 7458 748 7818 756
rect 6586 424 7258 426
rect 13297 424 13431 1290
rect 1805 402 7258 424
rect 1805 78 6648 402
rect 7052 78 7258 402
rect 1805 52 7258 78
rect 9144 386 25666 424
rect 9144 88 9188 386
rect 9462 332 25666 386
rect 9462 88 25447 332
rect 1805 46 6916 52
rect 9144 46 25447 88
rect 7456 -56 8966 -10
rect 7456 -262 7522 -56
rect 8864 -262 8966 -56
rect 7456 -302 8966 -262
<< via3 >>
rect 7532 808 8980 994
rect 7522 -262 8864 -56
<< metal4 >>
rect 1488 1136 2056 10916
rect 24592 1136 25160 6682
rect 1488 994 25160 1136
rect 1488 808 7532 994
rect 8980 808 25160 994
rect 1488 578 25160 808
rect 1488 568 24670 578
rect 7456 -28 8966 -10
rect 7456 -276 7518 -28
rect 8874 -276 8966 -28
rect 7456 -302 8966 -276
<< via4 >>
rect 7518 -56 8874 -28
rect 7518 -262 7522 -56
rect 7522 -262 8864 -56
rect 8864 -262 8874 -56
rect 7518 -276 8874 -262
<< metal5 >>
rect 789 46 1393 10802
rect 25314 7650 25904 9883
rect 25390 7316 25904 7650
rect 25314 46 25904 7316
rect 789 -28 25904 46
rect 789 -276 7518 -28
rect 8874 -276 25904 -28
rect 789 -507 25904 -276
rect 789 -558 25892 -507
use buffer_digital  buffer_digital_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 8708 0 1 68
box -274 0 415 576
use buffer_digital  buffer_digital_1
timestamp 1698771642
transform 1 0 7462 0 1 52
box -274 0 415 576
use charge_pump1_reverse  charge_pump1_reverse_0
timestamp 1698837094
transform 1 0 821 0 -1 27110
box -313 -3396 25321 25896
<< end >>
