magic
tech sky130A
magscale 1 2
timestamp 1698921260
<< pwell >>
rect 820 -8748 1040 -8700
rect 820 -8782 1146 -8748
<< poly >>
rect 148148 562 148246 1124
rect 148150 238 148248 344
rect 148150 136 148170 238
rect 148230 136 148248 238
rect 148150 110 148248 136
<< polycont >>
rect 148170 136 148230 238
<< locali >>
rect 148150 238 148244 254
rect 148150 136 148170 238
rect 148230 136 148244 238
rect 148150 110 148244 136
rect 820 -8714 1040 -8700
rect 820 -8766 840 -8714
rect 1012 -8748 1040 -8714
rect 1012 -8766 1146 -8748
rect 820 -8782 1146 -8766
rect 1206 -8784 1366 -8750
<< viali >>
rect 148170 136 148230 238
rect 840 -8766 1012 -8714
<< metal1 >>
rect -3767 48070 651 48072
rect -6574 47862 651 48070
rect -6574 46716 -3222 47862
rect -3782 -2028 -3222 46716
rect -3782 -5352 -3614 -2028
rect -3246 -5352 -3222 -2028
rect -3782 -48482 -3222 -5352
rect -3052 46572 -2492 46574
rect -3052 46544 440 46572
rect -3052 -6518 -2492 46544
rect -3052 -7226 -2964 -6518
rect -2554 -7226 -2492 -6518
rect -3052 -7300 -2492 -7226
rect -2380 44396 -1820 44402
rect -2380 44368 750 44396
rect -2380 44230 -1820 44368
rect -2380 42908 -2286 44230
rect -1922 42908 -1820 44230
rect -3052 -8660 -2492 -8508
rect -3052 -9368 -2964 -8660
rect -2554 -9368 -2492 -8660
rect -3052 -47164 -2492 -9368
rect -2380 -44988 -1820 42908
rect -1702 43308 -1142 43316
rect -1702 43280 804 43308
rect -1702 42834 -1142 43280
rect -1693 41992 -1142 42834
rect -1693 41586 -1588 41992
rect -1702 40534 -1588 41586
rect -1224 40534 -1142 41992
rect -1016 41744 -474 41752
rect -1016 41740 308 41744
rect -1702 -43900 -1142 40534
rect -1034 41716 308 41740
rect -1034 39544 -474 41716
rect -1034 38202 -1026 39544
rect -526 38202 -474 39544
rect -1034 -42336 -474 38202
rect -352 -41762 208 41136
rect 8730 4374 9252 4388
rect 8660 4316 9252 4374
rect 10397 4352 10537 4358
rect 10388 4346 10552 4352
rect 8660 3350 8916 4316
rect 10290 4182 10552 4346
rect 8606 3276 8962 3350
rect 8606 2824 8662 3276
rect 8896 2824 8962 3276
rect 8606 2784 8962 2824
rect 8730 2782 8802 2784
rect 896 938 1113 980
rect 10100 875 10226 3496
rect 10388 2256 10552 4182
rect 10966 3633 11060 3636
rect 14726 3633 14812 3636
rect 10965 3620 14819 3633
rect 10965 3599 10982 3620
rect 10966 3224 10982 3599
rect 11052 3612 14819 3620
rect 11052 3599 14738 3612
rect 11052 3224 11060 3599
rect 10966 3212 11060 3224
rect 14726 2858 14738 3599
rect 14798 3599 14819 3612
rect 14798 2858 14812 3599
rect 14726 2846 14812 2858
rect 10346 2186 10626 2256
rect 10346 1902 10408 2186
rect 10572 1902 10626 2186
rect 10346 1848 10626 1902
rect 151208 1850 151548 1882
rect 151208 1688 151236 1850
rect 151514 1688 151548 1850
rect 151208 1574 151548 1688
rect 9640 838 10226 875
rect 10100 836 10226 838
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 141714 440 143268 508
rect 148100 496 148136 1242
rect 148264 1160 148394 1168
rect 148264 1138 148320 1160
rect 148254 1108 148320 1138
rect 148384 1108 148394 1160
rect 148254 1104 148394 1108
rect 148264 1098 148394 1104
rect 148264 1096 148346 1098
rect 141923 -176 142237 440
rect 148259 384 148298 543
rect 148257 345 148437 384
rect 148150 238 148244 254
rect 148150 136 148170 238
rect 148230 136 148244 238
rect 148150 110 148244 136
rect 9349 -242 14172 -236
rect 9349 -264 14792 -242
rect 9349 -294 14078 -264
rect 9151 -335 14078 -294
rect 9349 -382 14078 -335
rect 14758 -382 14792 -264
rect 9349 -394 14792 -382
rect 9349 -402 14172 -394
rect 15072 -490 147551 -176
rect 148398 -2319 148437 345
rect 151372 382 151468 388
rect 151372 308 151384 382
rect 151456 308 151468 382
rect 151372 296 151468 308
rect 153290 366 153432 394
rect 150720 174 151114 214
rect 150720 68 150748 174
rect 151082 68 151114 174
rect 150720 46 151114 68
rect 151950 -83 152126 -74
rect 151950 -90 152127 -83
rect 151950 -158 151964 -90
rect 152116 -158 152127 -90
rect 151950 -170 152127 -158
rect 152073 -690 152127 -170
rect 152790 -782 152940 192
rect 153290 120 153310 366
rect 153414 120 153432 366
rect 153290 100 153432 120
rect 148384 -2336 154888 -2319
rect 148384 -2375 154901 -2336
rect 148384 -2535 154888 -2375
rect 148384 -2736 154896 -2535
rect 10780 -2892 10848 -2874
rect 10780 -3454 10786 -2892
rect 10457 -3484 10786 -3454
rect 10844 -3454 10848 -2892
rect 148400 -2952 154896 -2736
rect 10844 -3455 14406 -3454
rect 14458 -3455 14538 -3454
rect 10844 -3484 14727 -3455
rect 10457 -3489 14472 -3484
rect 10457 -3764 14406 -3489
rect 1612 -5797 3583 -5471
rect 1612 -7626 1938 -5797
rect 10457 -6583 10767 -3764
rect 14458 -4228 14472 -3489
rect 14524 -3489 14727 -3484
rect 14524 -4228 14538 -3489
rect 14458 -4242 14538 -4228
rect 14466 -4244 14516 -4242
rect 10994 -5486 11342 -5446
rect 10994 -5800 11040 -5486
rect 11300 -5800 11342 -5486
rect 10994 -5834 11342 -5800
rect 9611 -6645 10767 -6583
rect 9611 -6649 10697 -6645
rect 11057 -7675 11091 -5834
rect 820 -8714 1040 -8700
rect 820 -8766 840 -8714
rect 1012 -8766 1040 -8714
rect 820 -8782 1040 -8766
rect 1270 -8726 1432 -8714
rect 1270 -8780 1282 -8726
rect 1420 -8750 1432 -8726
rect 1420 -8780 1434 -8750
rect 1270 -8784 1434 -8780
rect 1650 -8919 1976 -8174
rect 1650 -9245 2969 -8919
rect 8486 -9204 9846 -9092
rect 11049 -9204 11121 -8826
rect 8486 -9214 11121 -9204
rect 1650 -9617 1976 -9245
rect 497 -9682 1976 -9617
rect 497 -9892 526 -9682
rect 1804 -9892 1976 -9682
rect 8486 -9776 8602 -9214
rect 9778 -9276 11121 -9214
rect 9778 -9776 9846 -9276
rect 8486 -9846 9846 -9776
rect 497 -9943 1976 -9892
rect -1034 -42364 -118 -42336
rect -1034 -42392 -474 -42364
rect -1702 -43916 384 -43900
rect -1698 -43928 384 -43916
rect -2380 -45006 324 -44988
rect -2360 -45016 324 -45006
rect -3052 -47190 184 -47164
rect -2908 -47192 184 -47190
rect -3782 -48692 545 -48482
<< via1 >>
rect -3614 -5352 -3246 -2028
rect -2964 -7226 -2554 -6518
rect -2286 42908 -1922 44230
rect -2964 -9368 -2554 -8660
rect -1588 40534 -1224 41992
rect -1026 38202 -526 39544
rect 8662 2824 8896 3276
rect 10982 3224 11052 3620
rect 14738 2858 14798 3612
rect 10408 1902 10572 2186
rect 151236 1688 151514 1850
rect 141758 508 143186 868
rect 148320 1108 148384 1160
rect 148170 136 148230 238
rect 14078 -382 14758 -264
rect 151384 308 151456 382
rect 150748 68 151082 174
rect 151964 -158 152116 -90
rect 153310 120 153414 366
rect 10786 -3484 10844 -2892
rect 14472 -4228 14524 -3484
rect 11040 -5800 11300 -5486
rect 840 -8766 1012 -8714
rect 1282 -8780 1420 -8726
rect 526 -9892 1804 -9682
rect 8602 -9776 9778 -9214
<< metal2 >>
rect 133308 87497 148018 87509
rect 133308 87428 148020 87497
rect 133308 87269 166338 87428
rect 146558 79019 166338 87269
rect -8551 44230 -1816 44386
rect -8551 42908 -2286 44230
rect -1922 42908 -1816 44230
rect -8551 42824 -1816 42908
rect -8468 41992 -1150 42074
rect -8468 40534 -1588 41992
rect -1224 40534 -1150 41992
rect -8468 40388 -1150 40534
rect -8260 39544 -494 39628
rect -8260 38202 -1026 39544
rect -526 38202 -494 39544
rect -8260 38108 -494 38202
rect -4264 4744 890 7690
rect 8568 6950 11198 7294
rect 8568 5410 8960 6950
rect 10878 5410 11198 6950
rect 8568 5070 11198 5410
rect -2626 3266 -1628 4744
rect 10674 3980 11034 5070
rect 10668 3636 11056 3980
rect 10668 3620 11060 3636
rect -2626 2398 -2468 3266
rect -1848 2398 -1628 3266
rect 8606 3276 8962 3350
rect 8606 2824 8662 3276
rect 8896 2824 8962 3276
rect 8606 2784 8962 2824
rect 10668 3224 10982 3620
rect 11052 3224 11060 3620
rect 10668 3212 11060 3224
rect 14726 3612 14812 3636
rect -2626 2132 -1628 2398
rect 10346 2186 10626 2256
rect 10346 1902 10408 2186
rect 10572 1902 10626 2186
rect 10346 1848 10626 1902
rect -5184 -680 674 1248
rect 1274 258 1688 260
rect 1156 234 1688 258
rect 1156 126 1198 234
rect 1600 126 1688 234
rect 1156 110 1688 126
rect 1156 108 1348 110
rect 1170 56 1630 58
rect 1156 34 1630 56
rect 1156 -54 1222 34
rect 1596 -54 1630 34
rect 1156 -94 1630 -54
rect -5108 -906 -4096 -680
rect 10668 -806 11056 3212
rect 14726 2858 14738 3612
rect 14798 2858 14812 3612
rect 15833 3272 16533 3315
rect 15833 3184 15888 3272
rect 16384 3184 16533 3272
rect 15833 3149 16533 3184
rect 148400 2983 148817 3023
rect 14726 2846 14812 2858
rect 148370 2667 154640 2983
rect 148370 2566 154648 2667
rect 148378 2250 154648 2566
rect 148383 1168 148425 2250
rect 151208 1850 151548 1882
rect 151208 1688 151236 1850
rect 151514 1688 151548 1850
rect 151208 1574 151548 1688
rect 148312 1160 148425 1168
rect 148312 1138 148320 1160
rect 148254 1108 148320 1138
rect 148384 1108 148425 1160
rect 148254 1104 148425 1108
rect 148312 1098 148425 1104
rect 148383 1097 148425 1098
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 141714 440 143268 508
rect 142442 156 142662 440
rect 151372 382 151468 390
rect 151372 308 151384 382
rect 151456 308 151468 382
rect 148148 238 148244 304
rect 12778 -64 147436 156
rect 148148 136 148170 238
rect 148230 142 148244 238
rect 150720 174 151114 214
rect 148230 136 148414 142
rect 148148 46 148414 136
rect 150720 68 150748 174
rect 151082 68 151114 174
rect 150720 46 151114 68
rect 151372 -74 151468 308
rect 153288 366 153436 396
rect 153288 120 153310 366
rect 153414 120 153436 366
rect 151372 -90 152128 -74
rect 151372 -158 151964 -90
rect 152116 -158 152128 -90
rect 151372 -170 152128 -158
rect 14046 -244 14792 -242
rect 153288 -244 153436 120
rect 14046 -264 153436 -244
rect 14046 -382 14078 -264
rect 14758 -382 153436 -264
rect 14046 -392 153436 -382
rect 14046 -394 14792 -392
rect 9786 -894 11056 -806
rect 12788 -808 150818 -588
rect -5108 -1554 -4990 -906
rect -4196 -1554 -4096 -906
rect -5108 -1672 -4096 -1554
rect -3754 -2028 -3176 -1728
rect -3754 -4654 -3614 -2028
rect -3766 -4766 -3614 -4654
rect -3778 -4966 -3614 -4766
rect -3754 -5352 -3614 -4966
rect -3246 -4654 -3176 -2028
rect -3246 -4966 9188 -4654
rect -3246 -5352 -3176 -4966
rect -3754 -5514 -3176 -5352
rect 8948 -5872 9188 -4966
rect 8948 -5920 9192 -5872
rect 8948 -6096 8982 -5920
rect 9160 -6096 9192 -5920
rect 8948 -6142 9192 -6096
rect 8948 -6150 9188 -6142
rect -3052 -6518 -2502 -6446
rect -3052 -7126 -2964 -6518
rect -3053 -7204 -2964 -7126
rect -3052 -7226 -2964 -7204
rect -2554 -7126 -2502 -6518
rect 10091 -6750 10344 -894
rect 150598 -1836 150818 -808
rect 152818 -1836 153038 -1276
rect 150598 -2056 153038 -1836
rect 10780 -2892 10848 -2874
rect 10780 -3484 10786 -2892
rect 10844 -3484 10848 -2892
rect 10780 -3494 10848 -3484
rect 14458 -3484 14538 -3454
rect 14458 -4228 14472 -3484
rect 14524 -4211 14538 -3484
rect 15850 -3792 16226 -3762
rect 15850 -3920 15898 -3792
rect 16176 -3920 16226 -3792
rect 15850 -3950 16226 -3920
rect 14524 -4228 14710 -4211
rect 14458 -4239 14710 -4228
rect 14458 -4242 14538 -4239
rect 14466 -4244 14516 -4242
rect 10994 -5486 11342 -5446
rect 10994 -5800 11040 -5486
rect 11300 -5800 11342 -5486
rect 10994 -5834 11342 -5800
rect -2554 -7204 2318 -7126
rect -2554 -7226 -2502 -7204
rect -3052 -7308 -2502 -7226
rect -3048 -8660 -2498 -8572
rect -3048 -8696 -2964 -8660
rect -3052 -8788 -2964 -8696
rect -3048 -9368 -2964 -8788
rect -2554 -8696 -2498 -8660
rect -2554 -8700 872 -8696
rect -2554 -8714 1040 -8700
rect -2554 -8766 840 -8714
rect 1012 -8766 1040 -8714
rect 1270 -8726 1432 -8714
rect 1270 -8750 1282 -8726
rect -2554 -8782 1040 -8766
rect 1206 -8780 1282 -8750
rect 1420 -8750 1432 -8726
rect 1420 -8780 2246 -8750
rect -2554 -8788 872 -8782
rect 1206 -8784 2246 -8780
rect -2554 -9368 -2498 -8788
rect -3048 -9434 -2498 -9368
rect 8486 -9214 9846 -9092
rect 420 -9682 1968 -9586
rect 420 -9704 526 -9682
rect -4326 -9892 526 -9704
rect 1804 -9892 1968 -9682
rect 8486 -9776 8602 -9214
rect 9778 -9776 9846 -9214
rect 8486 -9846 9846 -9776
rect -4326 -9940 1968 -9892
rect -4326 -12110 1058 -9940
rect 161022 -80316 166580 -79794
rect 147308 -87889 166580 -80316
rect 132474 -88070 166580 -87889
rect 132474 -88129 148006 -88070
rect 147370 -88143 148000 -88129
<< via2 >>
rect 8960 5410 10878 6950
rect -2468 2398 -1848 3266
rect 8662 2824 8896 3276
rect 10408 1902 10572 2186
rect 1198 126 1600 234
rect 1222 -54 1596 34
rect 15888 3184 16384 3272
rect 151236 1688 151514 1850
rect 141758 508 143186 868
rect 150748 68 151082 174
rect -4990 -1554 -4196 -906
rect 1606 -3340 2902 -2972
rect 8576 -3338 9764 -2976
rect 8982 -6096 9160 -5920
rect 10786 -3484 10844 -2892
rect 15898 -3920 16176 -3792
rect 11040 -5800 11300 -5486
rect 526 -9892 1804 -9682
rect 8602 -9776 9778 -9214
<< metal3 >>
rect -8526 6950 11258 7274
rect -8526 5410 8960 6950
rect 10878 5410 11258 6950
rect -8526 5070 11258 5410
rect -5176 3446 -2824 3456
rect -5176 3444 -824 3446
rect -5178 3266 -824 3444
rect -5178 3222 -2468 3266
rect -5178 2274 -4942 3222
rect -3104 2398 -2468 3222
rect -1848 2398 -824 3266
rect 8606 3276 8962 3350
rect 8606 2824 8662 3276
rect 8896 2824 8962 3276
rect 8606 2784 8962 2824
rect -3104 2276 -824 2398
rect -3104 2274 706 2276
rect -5178 1392 706 2274
rect 10346 2186 10626 2256
rect 10346 1902 10408 2186
rect 10572 1902 10626 2186
rect 10346 1848 10626 1902
rect -4218 1384 -824 1392
rect -6585 888 948 1054
rect 5229 802 5841 876
rect -6570 522 1696 591
rect -6582 392 1696 454
rect -6582 329 1699 392
rect -6584 258 1138 264
rect 1274 260 1390 264
rect 1274 258 1688 260
rect -6584 234 1688 258
rect -6584 136 1198 234
rect 1070 126 1198 136
rect 1600 126 1688 234
rect 1070 110 1688 126
rect 1088 48 1222 50
rect 1088 36 1630 48
rect -6575 34 1630 36
rect -6575 -54 1222 34
rect 1596 -54 1630 34
rect -6575 -94 1630 -54
rect -6575 -98 1222 -94
rect 10564 -375 10828 -374
rect 9549 -450 10851 -375
rect -5104 -906 780 -784
rect -5104 -1554 -4990 -906
rect -4196 -1554 780 -906
rect -5104 -1668 780 -1554
rect -104 -2878 780 -1668
rect -104 -2896 2032 -2878
rect -104 -2972 3252 -2896
rect -104 -3340 1606 -2972
rect 2902 -3340 3252 -2972
rect -104 -3454 3252 -3340
rect 8492 -2976 9900 -2888
rect 8492 -3338 8576 -2976
rect 9764 -3338 9900 -2976
rect 8492 -3448 9900 -3338
rect 10564 -2892 10851 -450
rect 10564 -3484 10786 -2892
rect 10844 -3484 10851 -2892
rect 8948 -5920 9192 -5872
rect 8948 -6096 8982 -5920
rect 9160 -6096 9192 -5920
rect 8948 -6142 9192 -6096
rect 8486 -9214 9846 -9092
rect 420 -9682 1968 -9586
rect 420 -9892 526 -9682
rect 1804 -9892 1968 -9682
rect 8486 -9776 8602 -9214
rect 9778 -9776 9846 -9214
rect 8486 -9846 9846 -9776
rect 420 -9940 1968 -9892
rect 10564 -10166 10851 -3484
rect 10994 -5486 11342 -5446
rect 10994 -5800 11040 -5486
rect 11300 -5800 11342 -5486
rect 10994 -5834 11342 -5800
rect -11674 -11775 10851 -10166
rect -11674 -11810 10710 -11775
rect 9785 -30482 11338 -30481
rect 11530 -30482 12425 30261
rect 15833 3272 16452 3314
rect 15833 3184 15888 3272
rect 16384 3184 16452 3272
rect 15833 3149 16452 3184
rect 151208 1850 151548 1882
rect 151208 1688 151236 1850
rect 151514 1688 151548 1850
rect 151208 1574 151548 1688
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 141714 440 143268 508
rect 142650 232 143030 440
rect 142650 174 151159 232
rect 142650 68 150748 174
rect 151082 68 151159 174
rect 142650 50 151159 68
rect 142650 -140 143030 50
rect 15062 -520 147620 -140
rect 142551 -1206 144558 -1108
rect 151336 -1204 151438 -1014
rect 149920 -1206 151438 -1204
rect 142264 -1210 151438 -1206
rect 142264 -1410 142634 -1210
rect 144396 -1310 151438 -1210
rect 144396 -1410 151378 -1310
rect 142264 -1502 151378 -1410
rect 15850 -3792 16226 -3762
rect 15850 -3824 15898 -3792
rect 15755 -3885 15898 -3824
rect 15850 -3920 15898 -3885
rect 16176 -3920 16226 -3792
rect 15850 -3950 16226 -3920
rect 9785 -31539 12425 -30482
rect 9785 -33235 10843 -31539
rect -12084 -95510 10770 -87288
<< via3 >>
rect -4942 2274 -3104 3222
rect -2468 2398 -1848 3266
rect 8662 2824 8896 3276
rect 10408 1902 10572 2186
rect -4990 -1554 -4196 -906
rect 8576 -3338 9764 -2976
rect 526 -9892 1804 -9682
rect 8602 -9776 9778 -9214
rect 11040 -5800 11300 -5486
rect 151236 1688 151514 1850
rect 141758 508 143186 868
rect 142634 -1410 144396 -1210
<< metal4 >>
rect -30725 103024 17476 108254
rect -30725 98072 17648 103024
rect 16921 94385 17619 98072
rect -4264 4744 890 7690
rect -5176 3222 -2824 3456
rect -5176 2274 -4942 3222
rect -3104 2274 -2824 3222
rect -5176 2076 -2824 2274
rect -2626 3266 -1628 4744
rect -2626 2398 -2468 3266
rect -1848 2398 -1628 3266
rect 8606 3278 8962 3350
rect 8606 2824 8654 3278
rect 8910 2824 8962 3278
rect 8606 2784 8962 2824
rect -2626 2132 -1628 2398
rect 9102 2186 11338 2252
rect 9102 1902 10408 2186
rect 10572 1902 11338 2186
rect 9102 1844 11338 1902
rect -5190 -682 1060 1212
rect 10930 128 11338 1844
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 141714 440 143268 508
rect 140356 128 141376 178
rect -5108 -906 -4096 -682
rect -5108 -1554 -4990 -906
rect -4196 -1554 -4096 -906
rect -5108 -1672 -4096 -1554
rect 10930 -866 141618 128
rect 8492 -2976 9900 -2888
rect -10346 -4062 -4938 -3018
rect 8492 -3338 8576 -2976
rect 9764 -3338 9900 -2976
rect 8492 -3448 9900 -3338
rect 10930 -4062 11338 -866
rect 140268 -870 141376 -866
rect 140268 -1102 141272 -870
rect 140268 -1210 144598 -1102
rect 140268 -1410 142634 -1210
rect 144396 -1410 144598 -1210
rect 140268 -1492 144598 -1410
rect -10346 -4470 11338 -4062
rect -10346 -4950 -4938 -4470
rect 10930 -5432 11338 -4470
rect 8528 -5486 11338 -5432
rect 8528 -5800 11040 -5486
rect 11300 -5800 11338 -5486
rect 8528 -5840 11338 -5800
rect 145536 -7134 146104 4496
rect 151204 1850 151550 1879
rect 151204 1688 151236 1850
rect 151514 1688 151550 1850
rect 151204 -700 151550 1688
rect 8486 -9214 9846 -9092
rect 420 -9682 1968 -9586
rect 420 -9704 526 -9682
rect -4326 -9892 526 -9704
rect 1804 -9892 1968 -9682
rect 8486 -9776 8602 -9214
rect 9778 -9776 9846 -9214
rect 8486 -9846 9846 -9776
rect -4326 -9940 1968 -9892
rect -4326 -12110 1058 -9940
<< via4 >>
rect -4942 2274 -3104 3222
rect -2468 2398 -1848 3266
rect 8654 3276 8910 3278
rect 8654 2824 8662 3276
rect 8662 2824 8896 3276
rect 8896 2824 8910 3276
rect 141758 508 143186 868
rect 8576 -3338 9764 -2976
rect 8602 -9776 9778 -9214
<< metal5 >>
rect 146169 5724 146682 5849
rect -10599 3278 9858 3463
rect -10599 3266 8654 3278
rect -10599 3222 -2468 3266
rect -10599 2274 -4942 3222
rect -3104 2398 -2468 3222
rect -1848 2824 8654 3266
rect 8910 2824 9858 3278
rect -1848 2398 9858 2824
rect -3104 2274 9858 2398
rect -10599 2088 9858 2274
rect 8483 -2702 9858 2088
rect 141714 944 143268 950
rect 138862 868 143292 944
rect 138862 508 141758 868
rect 143186 508 143292 868
rect 138862 442 143292 508
rect 13033 82 13831 297
rect 138874 82 140192 442
rect 141714 440 143268 442
rect 13033 -786 141618 82
rect 8480 -2726 9860 -2702
rect 13033 -2726 13831 -786
rect 138874 -852 140192 -786
rect 8458 -2976 13866 -2726
rect 8458 -3338 8576 -2976
rect 9764 -3338 13866 -2976
rect 8458 -3524 13866 -3338
rect 8480 -9214 9860 -3524
rect 146169 -7895 146759 5724
rect 8480 -9776 8602 -9214
rect 9778 -9776 9860 -9214
rect 8480 -10294 9860 -9776
rect 14840 -39909 15129 -39191
rect 15603 -98230 16321 -97802
rect -12568 -111168 16452 -98230
use cmfb_pmos  cmfb_pmos_0 ~/layout_files/differential_amplifier
timestamp 1698902756
transform 1 0 148450 0 1 -716
box -158 762 4965 2374
use comparator_final_compact  comparator_final_compact_0 ~/layout_files/differential_amplifier
timestamp 1698914177
transform -1 0 8641 0 1 -7048
box -2532 -2214 8653 1614
use full_stage_compact  full_stage_compact_0 ~/layout_files/differential_amplifier
timestamp 1698914652
transform 1 0 5194 0 1 -2632
box -4134 -770 6100 4979
use reconfigurable_CP  reconfigurable_CP_0
timestamp 1698913416
transform 1 0 16242 0 -1 63194
box -16084 -34774 130792 62844
use reconfigurable_CP  reconfigurable_CP_1
timestamp 1698913416
transform 1 0 15920 0 1 -63814
box -16084 -34774 130792 62844
use reference0_9  reference0_9_0
timestamp 1698902493
transform 0 -1 151950 1 0 -1574
box -66 -1120 1022 620
use reference  reference_0 ~/layout_files/differential_amplifier
timestamp 1698913862
transform 0 1 9942 -1 0 4408
box -32 -858 1956 500
use sky130_fd_pr__nfet_01v8_8Q9BPT  sky130_fd_pr__nfet_01v8_8Q9BPT_0
timestamp 1698902186
transform 1 0 148196 0 1 1206
box -108 -126 108 126
use sky130_fd_pr__nfet_01v8_V6PAVL  sky130_fd_pr__nfet_01v8_V6PAVL_0
timestamp 1698902186
transform 1 0 148198 0 1 446
box -108 -126 108 126
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/sky_pdk/sky130/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 1314 0 -1 -8528
box -38 -48 314 592
use source_follower_buffer  source_follower_buffer_0
timestamp 1698765072
transform 1 0 14893 0 1 -4323
box -217 -59 950 1017
use source_follower_buffer  source_follower_buffer_1
timestamp 1698765072
transform 1 0 14975 0 1 2765
box -217 -59 950 1017
<< labels >>
flabel metal5 15603 -105367 15617 -105363 0 FreeSans 4800 90 0 0 digital_gnd
flabel metal4 16921 102321 17619 103019 0 FreeSans 4800 90 0 0 digital_vdd
rlabel metal3 1158 358 1158 358 1 source
flabel space 8228 39660 9060 39802 0 FreeSans 3200 0 0 0 scan_out
flabel space 148376 1942 148438 2082 0 FreeSans 2400 90 0 0 vd1
flabel space 148306 -658 148460 -292 0 FreeSans 2400 90 0 0 vd2
flabel metal4 -30725 98072 -20543 108254 0 FreeSans 16000 0 0 0 digital_vdd_1.8V
flabel space -6158 -95630 2366 -87288 0 FreeSans 16000 0 0 0 clock(internal)_50MHz
flabel metal5 -6522 -108146 -1140 -101858 0 FreeSans 16000 0 0 0 Digital_gnd
flabel metal2 157929 79019 166338 87428 0 FreeSans 16000 0 0 0 vout+
flabel metal2 153340 2296 153890 2902 0 FreeSans 8000 0 0 0 vd1
flabel space 153456 -2960 154006 -2354 0 FreeSans 8000 0 0 0 vd2
flabel space 153424 -88070 161700 -79794 0 FreeSans 16000 0 0 0 vout-
flabel space -6574 46716 -5648 48142 0 FreeSans 8000 0 0 0 clk_external
flabel metal2 -7251 42824 -5689 44386 0 FreeSans 8000 0 0 0 scan_in
flabel metal2 -8468 40388 -6658 42012 0 FreeSans 8000 0 0 0 scan_en
flabel metal2 -8260 38108 -6042 39556 0 FreeSans 8000 0 0 0 reset
flabel space -5816 -100 -5606 34 0 FreeSans 1600 0 0 0 drain1
flabel space -5822 136 -5612 270 0 FreeSans 1600 0 0 0 drain2
rlabel metal3 1220 550 1220 550 1 ib1
rlabel metal1 912 962 912 962 1 ib2
rlabel space -5788 314 -5664 458 1 source
flabel space -5792 310 -5656 472 0 FreeSans 1600 0 0 0 source
flabel space -5886 612 -5706 680 0 FreeSans 1600 0 0 0 ib1
flabel space -5812 1068 -5638 1152 0 FreeSans 1600 0 0 0 ib2_1uA
flabel space -11610 -11898 -9966 -10254 0 FreeSans 8000 0 0 0 v_int-
flabel metal3 -8526 5070 -6322 7274 0 FreeSans 8000 0 0 0 v_int+
flabel metal4 -10346 -4950 -8000 -3018 0 FreeSans 6400 0 0 0 analog_vdd_1.8V
flabel space -10456 2110 -8262 3522 0 FreeSans 6400 0 0 0 analog_gnd
<< end >>
