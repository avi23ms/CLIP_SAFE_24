magic
tech sky130A
magscale 1 2
timestamp 1698684236
<< error_p >>
rect 94000 24654 94013 24670
rect 93972 24626 94013 24642
rect 44864 24546 44877 24562
rect 44836 24518 44877 24534
rect 89203 24498 90293 24506
rect 90361 24500 91393 24506
rect 89233 24490 89279 24498
rect 89329 24490 89375 24498
rect 89425 24490 89471 24498
rect 89521 24490 89567 24498
rect 89617 24490 89663 24498
rect 89713 24490 89759 24498
rect 89809 24490 89855 24498
rect 89905 24490 89951 24498
rect 90001 24490 90047 24498
rect 90097 24490 90143 24498
rect 90193 24490 90239 24498
rect 89175 24470 90321 24478
rect 90333 24472 91421 24478
rect 89205 24462 90267 24470
rect 89249 24418 90199 24420
rect 40067 24390 41157 24398
rect 41225 24392 42257 24398
rect 89277 24390 90171 24392
rect 40097 24382 40143 24390
rect 40193 24382 40239 24390
rect 40289 24382 40335 24390
rect 40385 24382 40431 24390
rect 40481 24382 40527 24390
rect 40577 24382 40623 24390
rect 40673 24382 40719 24390
rect 40769 24382 40815 24390
rect 40865 24382 40911 24390
rect 40961 24382 41007 24390
rect 41057 24382 41103 24390
rect 40039 24362 41185 24370
rect 41197 24364 42285 24370
rect 40069 24354 41131 24362
rect 40113 24310 41063 24312
rect 40141 24282 41035 24284
rect 89185 22712 90281 22716
rect 89487 22710 90281 22712
rect 89701 22708 90281 22710
rect 40049 22604 41145 22608
rect 40351 22602 41145 22604
rect 40565 22600 41145 22602
rect 76478 22324 76528 22326
rect 76574 22324 76624 22326
rect 76670 22324 76720 22326
rect 76766 22324 76816 22326
rect 76862 22324 76912 22326
rect 76958 22324 77008 22326
rect 77054 22324 77104 22326
rect 77150 22324 77200 22326
rect 77246 22324 77296 22326
rect 77342 22324 77392 22326
rect 77438 22324 77488 22326
rect 77534 22324 77584 22326
rect 77630 22324 77680 22326
rect 77726 22324 77776 22326
rect 77822 22324 77872 22326
rect 77918 22324 77968 22326
rect 78014 22324 78064 22326
rect 78110 22324 78160 22326
rect 78206 22324 78256 22326
rect 27246 22216 27296 22218
rect 27342 22216 27392 22218
rect 27438 22216 27488 22218
rect 27534 22216 27584 22218
rect 27630 22216 27680 22218
rect 27726 22216 27776 22218
rect 27822 22216 27872 22218
rect 27918 22216 27968 22218
rect 28014 22216 28064 22218
rect 28110 22216 28160 22218
rect 28206 22216 28256 22218
rect 28302 22216 28352 22218
rect 28398 22216 28448 22218
rect 28494 22216 28544 22218
rect 28590 22216 28640 22218
rect 28686 22216 28736 22218
rect 28782 22216 28832 22218
rect 28878 22216 28928 22218
rect 28974 22216 29024 22218
rect 29070 22216 29120 22218
rect 89207 20628 90303 20630
rect 89484 20626 90303 20628
rect 89698 20624 90303 20626
rect 82019 20608 83115 20612
rect 82019 20606 82828 20608
rect 82019 20604 82614 20606
rect 40071 20520 41167 20522
rect 40348 20518 41167 20520
rect 40562 20516 41167 20518
rect 32883 20500 33979 20504
rect 32883 20498 33692 20500
rect 32883 20496 33478 20498
rect 82019 18524 83115 18526
rect 82019 18522 82816 18524
rect 82019 18520 82602 18522
rect 40135 18434 41231 18438
rect 40370 18432 41231 18434
rect 40584 18430 41231 18432
rect 82029 16438 83125 16440
rect 82029 16436 82816 16438
rect 82029 16434 82602 16436
rect 40648 16346 41271 16348
rect 82037 14352 83133 14354
rect 82037 14350 82826 14352
rect 82037 14348 82612 14350
rect 82033 12266 83129 12270
rect 82033 12264 82834 12266
rect 82033 12262 82620 12264
rect 40143 12150 41239 12152
rect 40418 12148 41239 12150
rect 40632 12146 41239 12148
rect 40151 10064 41247 10068
rect 40442 10062 41247 10064
rect 40656 10060 41247 10062
<< error_s >>
rect 76198 22324 76242 22338
rect 76382 22324 76432 22326
rect 27062 22216 27106 22230
rect 99817 19406 99818 19412
rect 99789 19378 99818 19384
rect 89280 18796 90272 18800
rect 89760 18794 90272 18796
rect 89974 18792 90226 18794
rect 32914 18670 33906 18672
rect 32914 18668 33426 18670
rect 32960 18666 33212 18668
rect 99809 17312 99810 17332
rect 99854 17312 99920 17332
rect 99781 17284 99810 17304
rect 99854 17284 99892 17304
rect 90038 16708 90290 16710
rect 32914 16584 33906 16586
rect 32914 16582 33426 16584
rect 32960 16580 33212 16582
rect 32924 14498 33916 14500
rect 32924 14496 33436 14498
rect 32970 14494 33222 14496
rect 23590 12992 23732 12998
rect 23776 12992 23777 12998
rect 23618 12964 23732 12970
rect 23776 12964 23805 12970
rect 89328 12512 90320 12514
rect 89808 12510 90320 12512
rect 90022 12508 90274 12510
rect 32932 12412 33924 12416
rect 32932 12410 33444 12412
rect 32978 12408 33230 12410
rect 99858 11030 99906 11040
rect 99858 11002 99878 11012
rect 50405 10906 50406 10928
rect 50450 10906 50630 10928
rect 50377 10878 50406 10900
rect 50450 10878 50602 10900
rect 89352 10426 90344 10430
rect 89832 10424 90344 10426
rect 90046 10422 90298 10424
rect 23604 8806 23713 8824
rect 23757 8806 23758 8824
rect 72732 8822 72849 8846
rect 72893 8822 72894 8846
rect 23632 8778 23713 8796
rect 23757 8778 23786 8796
rect 72760 8794 72849 8818
rect 72893 8794 72922 8818
<< metal1 >>
rect 51968 2462 53780 2536
rect 51968 2426 52066 2462
rect 26284 2369 26928 2378
rect 26276 2318 26928 2369
rect 26276 1862 26368 2318
rect 26858 1862 26928 2318
rect 26276 1808 26928 1862
rect 51962 2104 52066 2426
rect 53698 2104 53780 2462
rect 73914 2298 74228 3334
rect 99360 2624 100962 2656
rect 99356 2596 100962 2624
rect 75770 2490 75882 2498
rect 75662 2484 75982 2490
rect 75544 2426 77224 2484
rect 51962 2008 53780 2104
rect 26276 -580 26418 1808
rect 25357 -722 27077 -580
rect 51962 -646 52310 2008
rect 75544 1994 75628 2426
rect 77148 1994 77224 2426
rect 75544 1928 77224 1994
rect 99356 2166 99424 2596
rect 100888 2166 100962 2596
rect 99356 2106 100962 2166
rect 50292 -686 53464 -646
rect 75562 -650 75982 1928
rect 99356 -544 99866 2106
rect 26634 -724 27076 -722
rect 73316 -744 77564 -650
rect 97756 -742 100870 -544
rect 73427 -762 77564 -744
rect 99356 -750 99866 -742
rect 50630 -1026 50698 -952
rect 24616 -1092 25116 -1078
rect 24616 -1124 25298 -1092
rect 24616 -1500 24672 -1124
rect 25030 -1294 25298 -1124
rect 25662 -1110 26476 -1078
rect 27288 -1082 27678 -1076
rect 27090 -1110 27678 -1082
rect 25662 -1138 26502 -1110
rect 27288 -1134 27678 -1110
rect 25662 -1142 26476 -1138
rect 25342 -1190 25412 -1178
rect 25342 -1254 25348 -1190
rect 25402 -1254 25412 -1190
rect 25342 -1272 25412 -1254
rect 25562 -1190 25628 -1178
rect 25562 -1254 25568 -1190
rect 25622 -1254 25628 -1190
rect 25562 -1272 25628 -1254
rect 26686 -1184 26752 -1178
rect 26686 -1248 26692 -1184
rect 26746 -1248 26752 -1184
rect 26686 -1272 26752 -1248
rect 26906 -1184 26972 -1178
rect 26906 -1248 26912 -1184
rect 26966 -1248 26972 -1184
rect 26906 -1272 26972 -1248
rect 25030 -1500 25116 -1294
rect 24616 -1542 25116 -1500
rect 27288 -1468 27342 -1134
rect 27626 -1468 27678 -1134
rect 27288 -1532 27678 -1468
rect 49636 -1112 50146 -1038
rect 50630 -1060 52918 -1026
rect 53462 -1048 53674 -1046
rect 50630 -1088 52930 -1060
rect 53462 -1074 54004 -1048
rect 50630 -1094 52918 -1088
rect 53606 -1092 54004 -1074
rect 73618 -1088 73666 -1040
rect 73618 -1090 77124 -1088
rect 49636 -1504 49690 -1112
rect 50054 -1504 50146 -1112
rect 50310 -1142 50368 -1126
rect 50310 -1202 50314 -1142
rect 50366 -1202 50368 -1142
rect 50310 -1224 50368 -1202
rect 50528 -1142 50586 -1126
rect 50528 -1202 50532 -1142
rect 50584 -1202 50586 -1142
rect 50528 -1224 50586 -1202
rect 53066 -1128 53124 -1110
rect 53066 -1188 53068 -1128
rect 53120 -1188 53124 -1128
rect 53066 -1208 53124 -1188
rect 53152 -1210 53210 -1112
rect 53282 -1128 53340 -1108
rect 53282 -1188 53284 -1128
rect 53336 -1188 53340 -1128
rect 53282 -1206 53340 -1188
rect 49636 -1546 50146 -1504
rect 53606 -1486 53652 -1092
rect 53952 -1486 54004 -1092
rect 53606 -1532 54004 -1486
rect 72774 -1192 73128 -1102
rect 73644 -1122 77124 -1090
rect 73644 -1150 77150 -1122
rect 77700 -1136 78274 -1108
rect 77852 -1144 78274 -1136
rect 73644 -1156 77124 -1150
rect 72774 -1518 72802 -1192
rect 73084 -1518 73128 -1192
rect 73302 -1204 73362 -1184
rect 73302 -1264 73306 -1204
rect 73360 -1264 73362 -1204
rect 73302 -1288 73362 -1264
rect 73520 -1204 73580 -1186
rect 73520 -1264 73522 -1204
rect 73576 -1264 73580 -1204
rect 73520 -1290 73580 -1264
rect 77302 -1190 77362 -1172
rect 77302 -1250 77304 -1190
rect 77358 -1250 77362 -1190
rect 77302 -1276 77362 -1250
rect 77518 -1190 77578 -1172
rect 77518 -1250 77522 -1190
rect 77576 -1250 77578 -1190
rect 77518 -1276 77578 -1250
rect 72774 -1542 73128 -1518
rect 77852 -1500 77878 -1144
rect 78236 -1500 78274 -1144
rect 77852 -1538 78274 -1500
rect 97180 -1136 97520 -1092
rect 97180 -1508 97214 -1136
rect 97478 -1508 97520 -1136
rect 98074 -1112 100378 -1098
rect 101178 -1112 101442 -1110
rect 98074 -1140 100430 -1112
rect 101004 -1140 101442 -1112
rect 98074 -1154 100378 -1140
rect 101178 -1156 101442 -1140
rect 97756 -1194 97816 -1174
rect 97756 -1254 97758 -1194
rect 97814 -1254 97816 -1194
rect 97756 -1270 97816 -1254
rect 97972 -1194 98034 -1180
rect 97972 -1254 97976 -1194
rect 98030 -1254 98034 -1194
rect 97972 -1272 98034 -1254
rect 100606 -1194 100664 -1178
rect 100606 -1254 100610 -1194
rect 100662 -1254 100664 -1194
rect 100606 -1268 100664 -1254
rect 100824 -1194 100882 -1178
rect 100824 -1254 100828 -1194
rect 100824 -1272 100882 -1254
rect 97180 -1540 97520 -1508
rect 101178 -1482 101222 -1156
rect 101400 -1482 101442 -1156
rect 101178 -1536 101442 -1482
<< via1 >>
rect 26368 1862 26858 2318
rect 52066 2104 53698 2462
rect 75628 1994 77148 2426
rect 99424 2166 100888 2596
rect 24672 -1500 25030 -1124
rect 25348 -1254 25402 -1190
rect 25568 -1254 25622 -1190
rect 26692 -1248 26746 -1184
rect 26912 -1248 26966 -1184
rect 27342 -1468 27626 -1134
rect 49690 -1504 50054 -1112
rect 50314 -1202 50366 -1142
rect 50532 -1202 50584 -1142
rect 53068 -1188 53120 -1128
rect 53284 -1188 53336 -1128
rect 53652 -1486 53952 -1092
rect 72802 -1518 73084 -1192
rect 73306 -1264 73360 -1204
rect 73522 -1264 73576 -1204
rect 77304 -1250 77358 -1190
rect 77522 -1250 77576 -1190
rect 77878 -1500 78236 -1144
rect 97214 -1508 97478 -1136
rect 97758 -1254 97814 -1194
rect 97976 -1254 98030 -1194
rect 100610 -1254 100662 -1194
rect 100828 -1254 100882 -1194
rect 101222 -1482 101400 -1156
<< metal2 >>
rect 98257 25316 98423 25355
rect 98257 25288 98460 25316
rect 98487 25288 98653 25341
rect 48985 25189 49151 25203
rect 48851 24573 49151 25189
rect 98257 24731 98653 25288
rect 98257 24697 98574 24731
rect 98376 24676 98460 24697
rect 23746 23322 25976 23478
rect 48176 23360 50496 23428
rect 72858 23402 75172 23484
rect 97378 23444 99910 23572
rect 97382 21472 99776 21476
rect 72828 21438 72984 21440
rect 23635 21416 23795 21418
rect 23635 21406 23826 21416
rect 23635 21372 25974 21406
rect 23698 21322 25974 21372
rect 72828 21374 72992 21438
rect 23734 21250 25974 21322
rect 48182 21262 50502 21330
rect 72828 21296 75156 21374
rect 97382 21360 99926 21472
rect 97394 21358 99926 21360
rect 97438 21346 99926 21358
rect 72842 21292 75156 21296
rect 23734 21234 25964 21250
rect 23734 21202 25984 21234
rect 25776 21150 25984 21202
rect 97398 19384 99786 19392
rect 23782 19178 25860 19238
rect 48254 19172 50574 19240
rect 72828 19220 75142 19302
rect 97398 19276 99842 19384
rect 23842 17068 25920 17128
rect 48290 17086 50610 17154
rect 72838 17128 75152 17210
rect 97448 17188 99892 17304
rect 23676 14984 26010 15056
rect 48324 14996 50644 15064
rect 72818 15030 75132 15112
rect 97464 15102 99908 15218
rect 23618 12898 25952 12970
rect 48286 12902 50606 12970
rect 72806 12960 75120 13042
rect 97424 12992 99872 13132
rect 97410 11012 99858 11044
rect 23610 10898 23756 10972
rect 23610 10806 25982 10898
rect 48282 10832 50602 10900
rect 72792 10868 75106 10950
rect 97410 10934 99878 11012
rect 97410 10904 99858 10934
rect 23640 10804 25982 10806
rect 97462 8826 99922 8904
rect 23632 8724 25966 8796
rect 48300 8714 50620 8782
rect 72760 8736 75074 8818
rect 24223 6921 24517 7575
rect 73381 6931 73547 7683
rect 24223 6907 24389 6921
rect 73934 3334 74232 3341
rect 51968 2462 53780 2536
rect 26338 2318 26928 2378
rect 26338 1862 26368 2318
rect 26858 1862 26928 2318
rect 51968 2104 52066 2462
rect 53698 2104 53780 2462
rect 73914 2298 74232 3334
rect 99360 2596 100962 2656
rect 51968 2008 53780 2104
rect 26338 1808 26928 1862
rect 24616 -1092 25116 -1078
rect 24616 -1124 25298 -1092
rect 24616 -1500 24672 -1124
rect 25030 -1294 25298 -1124
rect 27288 -1134 27678 -1076
rect 25342 -1184 27068 -1178
rect 25342 -1190 26692 -1184
rect 25342 -1254 25348 -1190
rect 25402 -1254 25568 -1190
rect 25622 -1248 26692 -1190
rect 26746 -1248 26912 -1184
rect 26966 -1248 27068 -1184
rect 25622 -1254 27068 -1248
rect 25342 -1260 27068 -1254
rect 25342 -1272 25910 -1260
rect 25030 -1500 25116 -1294
rect 24616 -1542 25116 -1500
rect 25830 -2138 25910 -1272
rect 26294 -1272 27068 -1260
rect 26294 -2138 26374 -1272
rect 27288 -1468 27342 -1134
rect 27626 -1468 27678 -1134
rect 27288 -1532 27678 -1468
rect 49636 -1112 50146 -1038
rect 53606 -1092 54004 -1048
rect 49636 -1504 49690 -1112
rect 50054 -1504 50146 -1112
rect 53066 -1126 53124 -1110
rect 53282 -1126 53340 -1108
rect 50310 -1128 53456 -1126
rect 50310 -1142 53068 -1128
rect 50310 -1202 50314 -1142
rect 50366 -1202 50532 -1142
rect 50584 -1188 53068 -1142
rect 53120 -1188 53284 -1128
rect 53336 -1188 53456 -1128
rect 50584 -1202 53456 -1188
rect 50310 -1224 53456 -1202
rect 49636 -1546 50146 -1504
rect 51408 -1226 52036 -1224
rect 25830 -2218 26374 -2138
rect 51408 -2148 51528 -1226
rect 51928 -2148 52036 -1226
rect 53606 -1486 53652 -1092
rect 53952 -1486 54004 -1092
rect 53606 -1532 54004 -1486
rect 72774 -1192 73128 -1102
rect 72774 -1518 72802 -1192
rect 73084 -1518 73128 -1192
rect 73302 -1196 73362 -1184
rect 73520 -1196 73580 -1186
rect 73934 -1196 74232 2298
rect 75544 2426 77224 2484
rect 75544 1994 75628 2426
rect 77148 1994 77224 2426
rect 99360 2166 99424 2596
rect 100888 2166 100962 2596
rect 99360 2106 100962 2166
rect 75544 1928 77224 1994
rect 77852 -1144 78274 -1108
rect 75252 -1196 75912 -1186
rect 77302 -1190 77362 -1172
rect 77302 -1196 77304 -1190
rect 73302 -1204 77304 -1196
rect 73302 -1264 73306 -1204
rect 73360 -1264 73522 -1204
rect 73576 -1226 77304 -1204
rect 73576 -1264 75302 -1226
rect 73302 -1276 75302 -1264
rect 73302 -1288 73362 -1276
rect 73520 -1290 73580 -1276
rect 73934 -1280 74232 -1276
rect 72774 -1542 73128 -1518
rect 51408 -2238 52036 -2148
rect 75252 -2162 75302 -1276
rect 75854 -1250 77304 -1226
rect 77358 -1196 77362 -1190
rect 77518 -1190 77578 -1172
rect 77518 -1196 77522 -1190
rect 77358 -1250 77522 -1196
rect 77576 -1196 77578 -1190
rect 77576 -1250 77680 -1196
rect 75854 -1276 77680 -1250
rect 75854 -2162 75912 -1276
rect 77852 -1500 77878 -1144
rect 78236 -1500 78274 -1144
rect 77852 -1538 78274 -1500
rect 97180 -1136 97520 -1092
rect 97180 -1508 97214 -1136
rect 97478 -1508 97520 -1136
rect 101178 -1156 101442 -1110
rect 97756 -1194 97816 -1176
rect 97756 -1206 97758 -1194
rect 97750 -1254 97758 -1206
rect 97814 -1206 97816 -1194
rect 97974 -1194 98034 -1180
rect 97974 -1206 97976 -1194
rect 97814 -1254 97976 -1206
rect 98030 -1206 98034 -1194
rect 100606 -1194 100664 -1178
rect 98934 -1206 99478 -1204
rect 100606 -1206 100610 -1194
rect 98030 -1254 100610 -1206
rect 100662 -1206 100664 -1194
rect 100824 -1194 100882 -1178
rect 100824 -1206 100828 -1194
rect 100662 -1254 100828 -1206
rect 100882 -1254 101006 -1206
rect 97750 -1264 101006 -1254
rect 97750 -1272 98972 -1264
rect 97974 -1274 98034 -1272
rect 97180 -1540 97520 -1508
rect 75252 -2232 75912 -2162
rect 98934 -2178 98972 -1272
rect 99434 -1272 101006 -1264
rect 99434 -2178 99478 -1272
rect 101178 -1482 101222 -1156
rect 101400 -1482 101442 -1156
rect 101178 -1536 101442 -1482
rect 98934 -2228 99478 -2178
<< via2 >>
rect 26368 1862 26858 2318
rect 52066 2104 53698 2462
rect 24672 -1500 25030 -1124
rect 25910 -2138 26294 -1260
rect 27342 -1468 27626 -1134
rect 49690 -1504 50054 -1112
rect 51528 -2148 51928 -1226
rect 53652 -1486 53952 -1092
rect 72802 -1518 73084 -1192
rect 75628 1994 77148 2426
rect 99424 2166 100888 2596
rect 75302 -2162 75854 -1226
rect 77878 -1500 78236 -1144
rect 97214 -1508 97478 -1136
rect 98972 -2178 99434 -1264
rect 101222 -1482 101400 -1156
<< metal3 >>
rect 99360 2596 100962 2656
rect 51968 2462 53780 2536
rect 26284 2318 26928 2378
rect 26284 1862 26368 2318
rect 26858 1862 26928 2318
rect 51968 2104 52066 2462
rect 53698 2104 53780 2462
rect 51968 2008 53780 2104
rect 75544 2426 77224 2484
rect 75544 1994 75628 2426
rect 77148 1994 77224 2426
rect 99360 2166 99424 2596
rect 100888 2166 100962 2596
rect 99360 2106 100962 2166
rect 75544 1928 77224 1994
rect 26284 1808 26928 1862
rect 12504 -1354 12638 173
rect 24616 -1094 25116 -1078
rect 24616 -1124 25306 -1094
rect 24616 -1354 24672 -1124
rect 12492 -1500 24672 -1354
rect 25030 -1278 25306 -1124
rect 27288 -1134 27678 -1076
rect 25830 -1260 26374 -1180
rect 25030 -1500 25116 -1278
rect 12492 -1538 25116 -1500
rect 12492 -1545 12638 -1538
rect 24616 -1542 25116 -1538
rect 25830 -2138 25910 -1260
rect 26294 -2138 26374 -1260
rect 27288 -1468 27342 -1134
rect 27626 -1354 27678 -1134
rect 37078 -1354 37194 -1054
rect 49636 -1112 50146 -1038
rect 49636 -1354 49690 -1112
rect 27626 -1408 38196 -1354
rect 39144 -1408 49690 -1354
rect 27626 -1468 49690 -1408
rect 27288 -1504 49690 -1468
rect 50054 -1504 50146 -1112
rect 53606 -1092 54004 -1048
rect 27288 -1538 50146 -1504
rect 49636 -1546 50146 -1538
rect 51408 -1226 52036 -1132
rect 25830 -2218 26374 -2138
rect 51408 -2148 51528 -1226
rect 51928 -2148 52036 -1226
rect 53606 -1486 53652 -1092
rect 53952 -1354 54004 -1092
rect 61640 -1354 61774 179
rect 72774 -1192 73128 -1102
rect 77852 -1144 78274 -1108
rect 72774 -1354 72802 -1192
rect 53952 -1486 72802 -1354
rect 53606 -1518 72802 -1486
rect 73084 -1518 73128 -1192
rect 53606 -1538 73128 -1518
rect 72774 -1542 73128 -1538
rect 75252 -1226 75912 -1186
rect 51408 -2238 52036 -2148
rect 75252 -2162 75302 -1226
rect 75854 -2162 75912 -1226
rect 77852 -1500 77878 -1144
rect 78236 -1354 78274 -1144
rect 86182 -1354 86420 -954
rect 97180 -1136 97520 -1092
rect 97180 -1354 97214 -1136
rect 78236 -1500 97214 -1354
rect 77852 -1508 97214 -1500
rect 97478 -1508 97520 -1136
rect 101178 -1156 101442 -1110
rect 77852 -1538 97520 -1508
rect 86182 -1554 86420 -1538
rect 97180 -1540 97520 -1538
rect 98934 -1264 99478 -1204
rect 75252 -2232 75912 -2162
rect 98934 -2178 98972 -1264
rect 99434 -2178 99478 -1264
rect 101178 -1482 101222 -1156
rect 101400 -1354 101442 -1156
rect 111046 -1354 111180 341
rect 101400 -1482 111194 -1354
rect 101178 -1538 111194 -1482
rect 111046 -1551 111180 -1538
rect 98934 -2228 99478 -2178
<< via3 >>
rect 26368 1862 26858 2318
rect 52066 2104 53698 2462
rect 75628 1994 77148 2426
rect 99424 2166 100888 2596
rect 25910 -2138 26294 -1260
rect 51528 -2148 51928 -1226
rect 75302 -2162 75854 -1226
rect 98972 -2178 99434 -1264
<< metal4 >>
rect 24255 10342 25585 24461
rect 23804 9012 25801 10342
rect 48690 9442 49898 24074
rect 48394 8234 50364 9442
rect 97545 8026 99805 24444
rect 99360 2596 100962 2656
rect 51968 2462 53780 2536
rect 51968 2104 52066 2462
rect 53698 2104 53780 2462
rect 51968 2008 53780 2104
rect 75544 2426 77224 2484
rect 75544 1994 75628 2426
rect 77148 1994 77224 2426
rect 99360 2166 99424 2596
rect 100888 2166 100962 2596
rect 99360 2106 100962 2166
rect 75544 1928 77224 1994
rect 25830 -1260 26374 -1180
rect 25830 -2138 25910 -1260
rect 26294 -2138 26374 -1260
rect 25830 -2218 26374 -2138
rect 51408 -1226 52036 -1132
rect 51408 -2148 51528 -1226
rect 51928 -2148 52036 -1226
rect 51408 -2238 52036 -2148
rect 75252 -1226 75912 -1186
rect 75252 -2162 75302 -1226
rect 75854 -2162 75912 -1226
rect 75252 -2232 75912 -2162
rect 98934 -1264 99478 -1204
rect 98934 -2178 98972 -1264
rect 99434 -2178 99478 -1264
rect 98934 -2228 99478 -2178
<< via4 >>
rect 25910 -2138 26294 -1260
rect 51528 -2148 51928 -1226
rect 75302 -2162 75854 -1226
rect 98972 -2178 99434 -1264
<< metal5 >>
rect 56 -1622 660 8374
rect 25830 -1260 26374 -1180
rect 25830 -1622 25910 -1260
rect 56 -2138 25910 -1622
rect 26294 -1622 26374 -1260
rect 51408 -1226 52036 -1132
rect 51408 -1622 51528 -1226
rect 26294 -1664 37908 -1622
rect 39228 -1664 51528 -1622
rect 26294 -2138 51528 -1664
rect 56 -2148 51528 -2138
rect 51928 -1622 52036 -1226
rect 75230 -1226 75930 -1178
rect 75230 -1622 75302 -1226
rect 51928 -2148 75302 -1622
rect 56 -2162 75302 -2148
rect 75854 -1622 75930 -1226
rect 98934 -1264 99478 -1204
rect 98934 -1622 98972 -1264
rect 75854 -2162 98972 -1622
rect 56 -2178 98972 -2162
rect 99434 -1622 99478 -1264
rect 123063 -1622 123653 3937
rect 99434 -2178 123670 -1622
rect 56 -2226 123670 -2178
rect 51408 -2238 52036 -2226
rect 75230 -2246 75930 -2226
rect 98934 -2228 99478 -2226
use buffer_digital  buffer_digital_1 ~/Desktop/charge_pumps2/layout_files
timestamp 1698389822
transform 1 0 25360 0 1 -1292
box -274 0 412 576
use buffer_digital  buffer_digital_3
timestamp 1698389822
transform 1 0 26706 0 1 -1278
box -274 0 412 576
use buffer_digital  buffer_digital_4
timestamp 1698389822
transform 1 0 50324 0 1 -1242
box -274 0 412 576
use buffer_digital  buffer_digital_5
timestamp 1698389822
transform 1 0 53078 0 1 -1228
box -274 0 412 576
use buffer_digital  buffer_digital_6
timestamp 1698389822
transform 1 0 73316 0 1 -1304
box -274 0 412 576
use buffer_digital  buffer_digital_7
timestamp 1698389822
transform 1 0 77316 0 1 -1290
box -274 0 412 576
use buffer_digital  buffer_digital_8
timestamp 1698389822
transform 1 0 97770 0 1 -1294
box -274 0 412 576
use buffer_digital  buffer_digital_9
timestamp 1698389822
transform 1 0 100620 0 1 -1294
box -274 0 412 576
use charge_pump1  charge_pump1_0
timestamp 1698684236
transform 1 0 28 0 1 7576
box -313 -7588 25321 19132
use charge_pump1  charge_pump1_1
timestamp 1698684236
transform 1 0 49164 0 1 7592
box -313 -7588 25321 19132
use charge_pump1  charge_pump1_2
timestamp 1698684236
transform 1 0 98570 0 1 7716
box -313 -7588 25321 19132
use charge_pump2  charge_pump2_0
timestamp 1698684236
transform 1 0 24536 0 -1 24556
box -313 -3396 25321 25892
use charge_pump2  charge_pump2_1
timestamp 1698684236
transform 1 0 73672 0 -1 24664
box -313 -3396 25321 25892
<< end >>
