* SPICE3 file created from nmos_dnw.ext - technology: sky130A

X0 dw_n418_1130# a_590_1174# a_606_1858# dw_n418_1130# sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.13 ps=1.46 w=0.42 l=0.15
X1 a_200_1200# a_0_1172# dw_n418_1130# dw_n418_1130# sky130_fd_pr__nfet_01v8 ad=1.65 pd=7.1 as=1.65 ps=7.1 w=3 l=1
X2 dw_n418_1130# a_590_1174# a_480_1200# dw_n418_1130# sky130_fd_pr__nfet_01v8 ad=1.65 pd=7.1 as=1.65 ps=7.1 w=3 l=1
X3 a_110_1858# a_0_1172# dw_n418_1130# dw_n418_1130# sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.126 ps=1.44 w=0.42 l=0.15
C0 dw_n418_1130# VSUBS 7.81f **FLOATING
