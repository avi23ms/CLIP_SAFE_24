magic
tech sky130A
magscale 1 2
timestamp 1699103691
<< nwell >>
rect -401 188 401 226
rect -497 -226 497 188
<< pmos >>
rect -399 -126 -369 126
rect -303 -126 -273 126
rect -207 -126 -177 126
rect -111 -126 -81 126
rect -15 -126 15 126
rect 81 -126 111 126
rect 177 -126 207 126
rect 273 -126 303 126
rect 369 -126 399 126
<< pdiff >>
rect -461 114 -399 126
rect -461 -114 -449 114
rect -415 -114 -399 114
rect -461 -126 -399 -114
rect -369 114 -303 126
rect -369 -114 -353 114
rect -319 -114 -303 114
rect -369 -126 -303 -114
rect -273 114 -207 126
rect -273 -114 -257 114
rect -223 -114 -207 114
rect -273 -126 -207 -114
rect -177 114 -111 126
rect -177 -114 -161 114
rect -127 -114 -111 114
rect -177 -126 -111 -114
rect -81 114 -15 126
rect -81 -114 -65 114
rect -31 -114 -15 114
rect -81 -126 -15 -114
rect 15 114 81 126
rect 15 -114 31 114
rect 65 -114 81 114
rect 15 -126 81 -114
rect 111 114 177 126
rect 111 -114 127 114
rect 161 -114 177 114
rect 111 -126 177 -114
rect 207 114 273 126
rect 207 -114 223 114
rect 257 -114 273 114
rect 207 -126 273 -114
rect 303 114 369 126
rect 303 -114 319 114
rect 353 -114 369 114
rect 303 -126 369 -114
rect 399 114 461 126
rect 399 -114 415 114
rect 449 -114 461 114
rect 399 -126 461 -114
<< pdiffc >>
rect -449 -114 -415 114
rect -353 -114 -319 114
rect -257 -114 -223 114
rect -161 -114 -127 114
rect -65 -114 -31 114
rect 31 -114 65 114
rect 127 -114 161 114
rect 223 -114 257 114
rect 319 -114 353 114
rect 415 -114 449 114
<< poly >>
rect -321 207 -255 223
rect -321 173 -305 207
rect -271 173 -255 207
rect -321 157 -255 173
rect -129 207 -63 223
rect -129 173 -113 207
rect -79 173 -63 207
rect -129 157 -63 173
rect 63 207 129 223
rect 63 173 79 207
rect 113 173 129 207
rect 63 157 129 173
rect 255 207 321 223
rect 255 173 271 207
rect 305 173 321 207
rect 255 157 321 173
rect -399 126 -369 152
rect -303 126 -273 157
rect -207 126 -177 152
rect -111 126 -81 157
rect -15 126 15 152
rect 81 126 111 157
rect 177 126 207 152
rect 273 126 303 157
rect 369 126 399 152
rect -399 -157 -369 -126
rect -303 -152 -273 -126
rect -207 -157 -177 -126
rect -111 -152 -81 -126
rect -15 -157 15 -126
rect 81 -152 111 -126
rect 177 -157 207 -126
rect 273 -152 303 -126
rect 369 -157 399 -126
rect -417 -173 -351 -157
rect -417 -207 -401 -173
rect -367 -207 -351 -173
rect -417 -223 -351 -207
rect -225 -173 -159 -157
rect -225 -207 -209 -173
rect -175 -207 -159 -173
rect -225 -223 -159 -207
rect -33 -173 33 -157
rect -33 -207 -17 -173
rect 17 -207 33 -173
rect -33 -223 33 -207
rect 159 -173 225 -157
rect 159 -207 175 -173
rect 209 -207 225 -173
rect 159 -223 225 -207
rect 351 -173 417 -157
rect 351 -207 367 -173
rect 401 -207 417 -173
rect 351 -223 417 -207
<< polycont >>
rect -305 173 -271 207
rect -113 173 -79 207
rect 79 173 113 207
rect 271 173 305 207
rect -401 -207 -367 -173
rect -209 -207 -175 -173
rect -17 -207 17 -173
rect 175 -207 209 -173
rect 367 -207 401 -173
<< locali >>
rect -321 173 -305 207
rect -271 173 -255 207
rect -129 173 -113 207
rect -79 173 -63 207
rect 63 173 79 207
rect 113 173 129 207
rect 255 173 271 207
rect 305 173 321 207
rect -449 114 -415 130
rect -449 -130 -415 -114
rect -353 114 -319 130
rect -353 -130 -319 -114
rect -257 114 -223 130
rect -257 -130 -223 -114
rect -161 114 -127 130
rect -161 -130 -127 -114
rect -65 114 -31 130
rect -65 -130 -31 -114
rect 31 114 65 130
rect 31 -130 65 -114
rect 127 114 161 130
rect 127 -130 161 -114
rect 223 114 257 130
rect 223 -130 257 -114
rect 319 114 353 130
rect 319 -130 353 -114
rect 415 114 449 130
rect 415 -130 449 -114
rect -417 -207 -401 -173
rect -367 -207 -351 -173
rect -225 -207 -209 -173
rect -175 -207 -159 -173
rect -33 -207 -17 -173
rect 17 -207 33 -173
rect 159 -207 175 -173
rect 209 -207 225 -173
rect 351 -207 367 -173
rect 401 -207 417 -173
<< viali >>
rect -449 -114 -415 114
rect -353 -114 -319 114
rect -257 -114 -223 114
rect -161 -114 -127 114
rect -65 -114 -31 114
rect 31 -114 65 114
rect 127 -114 161 114
rect 223 -114 257 114
rect 319 -114 353 114
rect 415 -114 449 114
<< metal1 >>
rect -455 114 -409 126
rect -455 -114 -449 114
rect -415 -114 -409 114
rect -455 -126 -409 -114
rect -359 114 -313 126
rect -359 -114 -353 114
rect -319 -114 -313 114
rect -359 -126 -313 -114
rect -263 114 -217 126
rect -263 -114 -257 114
rect -223 -114 -217 114
rect -263 -126 -217 -114
rect -167 114 -121 126
rect -167 -114 -161 114
rect -127 -114 -121 114
rect -167 -126 -121 -114
rect -71 114 -25 126
rect -71 -114 -65 114
rect -31 -114 -25 114
rect -71 -126 -25 -114
rect 25 114 71 126
rect 25 -114 31 114
rect 65 -114 71 114
rect 25 -126 71 -114
rect 121 114 167 126
rect 121 -114 127 114
rect 161 -114 167 114
rect 121 -126 167 -114
rect 217 114 263 126
rect 217 -114 223 114
rect 257 -114 263 114
rect 217 -126 263 -114
rect 313 114 359 126
rect 313 -114 319 114
rect 353 -114 359 114
rect 313 -126 359 -114
rect 409 114 455 126
rect 409 -114 415 114
rect 449 -114 455 114
rect 409 -126 455 -114
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.26 l 0.15 m 1 nf 9 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
